module nv_ram_rwsp( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_clk, // @[:@6.4]
  input         io_re, // @[:@6.4]
  input         io_we, // @[:@6.4]
  input         io_ore, // @[:@6.4]
  input  [6:0]  io_ra, // @[:@6.4]
  input  [6:0]  io_wa, // @[:@6.4]
  input  [31:0] io_pwrbus_ram_pd, // @[:@6.4]
  input  [10:0] io_di, // @[:@6.4]
  output [10:0] io_dout // @[:@6.4]
);
  reg [10:0] mem_0; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_0;
  reg [10:0] mem_1; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_1;
  reg [10:0] mem_2; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_2;
  reg [10:0] mem_3; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_3;
  reg [10:0] mem_4; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_4;
  reg [10:0] mem_5; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_5;
  reg [10:0] mem_6; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_6;
  reg [10:0] mem_7; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_7;
  reg [10:0] mem_8; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_8;
  reg [10:0] mem_9; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_9;
  reg [10:0] mem_10; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_10;
  reg [10:0] mem_11; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_11;
  reg [10:0] mem_12; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_12;
  reg [10:0] mem_13; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_13;
  reg [10:0] mem_14; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_14;
  reg [10:0] mem_15; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_15;
  reg [10:0] mem_16; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_16;
  reg [10:0] mem_17; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_17;
  reg [10:0] mem_18; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_18;
  reg [10:0] mem_19; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_19;
  reg [10:0] mem_20; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_20;
  reg [10:0] mem_21; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_21;
  reg [10:0] mem_22; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_22;
  reg [10:0] mem_23; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_23;
  reg [10:0] mem_24; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_24;
  reg [10:0] mem_25; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_25;
  reg [10:0] mem_26; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_26;
  reg [10:0] mem_27; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_27;
  reg [10:0] mem_28; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_28;
  reg [10:0] mem_29; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_29;
  reg [10:0] mem_30; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_30;
  reg [10:0] mem_31; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_31;
  reg [10:0] mem_32; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_32;
  reg [10:0] mem_33; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_33;
  reg [10:0] mem_34; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_34;
  reg [10:0] mem_35; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_35;
  reg [10:0] mem_36; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_36;
  reg [10:0] mem_37; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_37;
  reg [10:0] mem_38; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_38;
  reg [10:0] mem_39; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_39;
  reg [10:0] mem_40; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_40;
  reg [10:0] mem_41; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_41;
  reg [10:0] mem_42; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_42;
  reg [10:0] mem_43; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_43;
  reg [10:0] mem_44; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_44;
  reg [10:0] mem_45; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_45;
  reg [10:0] mem_46; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_46;
  reg [10:0] mem_47; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_47;
  reg [10:0] mem_48; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_48;
  reg [10:0] mem_49; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_49;
  reg [10:0] mem_50; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_50;
  reg [10:0] mem_51; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_51;
  reg [10:0] mem_52; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_52;
  reg [10:0] mem_53; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_53;
  reg [10:0] mem_54; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_54;
  reg [10:0] mem_55; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_55;
  reg [10:0] mem_56; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_56;
  reg [10:0] mem_57; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_57;
  reg [10:0] mem_58; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_58;
  reg [10:0] mem_59; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_59;
  reg [10:0] mem_60; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_60;
  reg [10:0] mem_61; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_61;
  reg [10:0] mem_62; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_62;
  reg [10:0] mem_63; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_63;
  reg [10:0] mem_64; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_64;
  reg [10:0] mem_65; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_65;
  reg [10:0] mem_66; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_66;
  reg [10:0] mem_67; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_67;
  reg [10:0] mem_68; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_68;
  reg [10:0] mem_69; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_69;
  reg [10:0] mem_70; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_70;
  reg [10:0] mem_71; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_71;
  reg [10:0] mem_72; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_72;
  reg [10:0] mem_73; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_73;
  reg [10:0] mem_74; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_74;
  reg [10:0] mem_75; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_75;
  reg [10:0] mem_76; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_76;
  reg [10:0] mem_77; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_77;
  reg [10:0] mem_78; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_78;
  reg [10:0] mem_79; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_79;
  reg [10:0] mem_80; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_80;
  reg [10:0] mem_81; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_81;
  reg [10:0] mem_82; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_82;
  reg [10:0] mem_83; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_83;
  reg [10:0] mem_84; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_84;
  reg [10:0] mem_85; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_85;
  reg [10:0] mem_86; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_86;
  reg [10:0] mem_87; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_87;
  reg [10:0] mem_88; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_88;
  reg [10:0] mem_89; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_89;
  reg [10:0] mem_90; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_90;
  reg [10:0] mem_91; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_91;
  reg [10:0] mem_92; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_92;
  reg [10:0] mem_93; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_93;
  reg [10:0] mem_94; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_94;
  reg [10:0] mem_95; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_95;
  reg [10:0] mem_96; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_96;
  reg [10:0] mem_97; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_97;
  reg [10:0] mem_98; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_98;
  reg [10:0] mem_99; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_99;
  reg [10:0] mem_100; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_100;
  reg [10:0] mem_101; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_101;
  reg [10:0] mem_102; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_102;
  reg [10:0] mem_103; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_103;
  reg [10:0] mem_104; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_104;
  reg [10:0] mem_105; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_105;
  reg [10:0] mem_106; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_106;
  reg [10:0] mem_107; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_107;
  reg [10:0] mem_108; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_108;
  reg [10:0] mem_109; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_109;
  reg [10:0] mem_110; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_110;
  reg [10:0] mem_111; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_111;
  reg [10:0] mem_112; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_112;
  reg [10:0] mem_113; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_113;
  reg [10:0] mem_114; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_114;
  reg [10:0] mem_115; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_115;
  reg [10:0] mem_116; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_116;
  reg [10:0] mem_117; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_117;
  reg [10:0] mem_118; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_118;
  reg [10:0] mem_119; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_119;
  reg [10:0] mem_120; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_120;
  reg [10:0] mem_121; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_121;
  reg [10:0] mem_122; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_122;
  reg [10:0] mem_123; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_123;
  reg [10:0] mem_124; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_124;
  reg [10:0] mem_125; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_125;
  reg [10:0] mem_126; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_126;
  reg [10:0] mem_127; // @[nv_ram_rwsp.scala 32:18:@8.4]
  reg [31:0] _RAND_127;
  reg [6:0] ra_d; // @[nv_ram_rwsp.scala 33:19:@9.4]
  reg [31:0] _RAND_128;
  reg [10:0] dout_r; // @[nv_ram_rwsp.scala 34:21:@10.4]
  reg [31:0] _RAND_129;
  wire [10:0] _GEN_0; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_1; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_2; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_3; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_4; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_5; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_6; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_7; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_8; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_9; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_10; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_11; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_12; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_13; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_14; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_15; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_16; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_17; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_18; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_19; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_20; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_21; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_22; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_23; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_24; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_25; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_26; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_27; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_28; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_29; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_30; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_31; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_32; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_33; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_34; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_35; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_36; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_37; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_38; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_39; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_40; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_41; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_42; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_43; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_44; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_45; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_46; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_47; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_48; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_49; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_50; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_51; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_52; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_53; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_54; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_55; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_56; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_57; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_58; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_59; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_60; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_61; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_62; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_63; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_64; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_65; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_66; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_67; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_68; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_69; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_70; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_71; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_72; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_73; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_74; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_75; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_76; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_77; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_78; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_79; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_80; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_81; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_82; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_83; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_84; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_85; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_86; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_87; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_88; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_89; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_90; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_91; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_92; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_93; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_94; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_95; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_96; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_97; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_98; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_99; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_100; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_101; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_102; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_103; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_104; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_105; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_106; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_107; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_108; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_109; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_110; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_111; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_112; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_113; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_114; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_115; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_116; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_117; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_118; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_119; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_120; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_121; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_122; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_123; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_124; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_125; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_126; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_127; // @[nv_ram_rwsp.scala 37:20:@12.6]
  wire [10:0] _GEN_258; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_259; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_260; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_261; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_262; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_263; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_264; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_265; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_266; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_267; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_268; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_269; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_270; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_271; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_272; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_273; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_274; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_275; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_276; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_277; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_278; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_279; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_280; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_281; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_282; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_283; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_284; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_285; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_286; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_287; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_288; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_289; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_290; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_291; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_292; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_293; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_294; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_295; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_296; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_297; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_298; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_299; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_300; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_301; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_302; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_303; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_304; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_305; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_306; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_307; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_308; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_309; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_310; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_311; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_312; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_313; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_314; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_315; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_316; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_317; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_318; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_319; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_320; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_321; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_322; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_323; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_324; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_325; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_326; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_327; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_328; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_329; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_330; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_331; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_332; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_333; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_334; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_335; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_336; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_337; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_338; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_339; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_340; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_341; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_342; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_343; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_344; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_345; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_346; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_347; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_348; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_349; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_350; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_351; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_352; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_353; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_354; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_355; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_356; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_357; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_358; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_359; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_360; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_361; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_362; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_363; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_364; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_365; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_366; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_367; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_368; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_369; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_370; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_371; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_372; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_373; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_374; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_375; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_376; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_377; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_378; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_379; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_380; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_381; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_382; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_383; // @[nv_ram_rwsp.scala 44:16:@18.6]
  wire [10:0] _GEN_384; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_0 = 7'h0 == io_wa ? io_di : mem_0; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_1 = 7'h1 == io_wa ? io_di : mem_1; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_2 = 7'h2 == io_wa ? io_di : mem_2; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_3 = 7'h3 == io_wa ? io_di : mem_3; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_4 = 7'h4 == io_wa ? io_di : mem_4; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_5 = 7'h5 == io_wa ? io_di : mem_5; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_6 = 7'h6 == io_wa ? io_di : mem_6; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_7 = 7'h7 == io_wa ? io_di : mem_7; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_8 = 7'h8 == io_wa ? io_di : mem_8; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_9 = 7'h9 == io_wa ? io_di : mem_9; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_10 = 7'ha == io_wa ? io_di : mem_10; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_11 = 7'hb == io_wa ? io_di : mem_11; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_12 = 7'hc == io_wa ? io_di : mem_12; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_13 = 7'hd == io_wa ? io_di : mem_13; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_14 = 7'he == io_wa ? io_di : mem_14; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_15 = 7'hf == io_wa ? io_di : mem_15; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_16 = 7'h10 == io_wa ? io_di : mem_16; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_17 = 7'h11 == io_wa ? io_di : mem_17; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_18 = 7'h12 == io_wa ? io_di : mem_18; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_19 = 7'h13 == io_wa ? io_di : mem_19; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_20 = 7'h14 == io_wa ? io_di : mem_20; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_21 = 7'h15 == io_wa ? io_di : mem_21; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_22 = 7'h16 == io_wa ? io_di : mem_22; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_23 = 7'h17 == io_wa ? io_di : mem_23; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_24 = 7'h18 == io_wa ? io_di : mem_24; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_25 = 7'h19 == io_wa ? io_di : mem_25; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_26 = 7'h1a == io_wa ? io_di : mem_26; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_27 = 7'h1b == io_wa ? io_di : mem_27; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_28 = 7'h1c == io_wa ? io_di : mem_28; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_29 = 7'h1d == io_wa ? io_di : mem_29; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_30 = 7'h1e == io_wa ? io_di : mem_30; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_31 = 7'h1f == io_wa ? io_di : mem_31; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_32 = 7'h20 == io_wa ? io_di : mem_32; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_33 = 7'h21 == io_wa ? io_di : mem_33; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_34 = 7'h22 == io_wa ? io_di : mem_34; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_35 = 7'h23 == io_wa ? io_di : mem_35; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_36 = 7'h24 == io_wa ? io_di : mem_36; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_37 = 7'h25 == io_wa ? io_di : mem_37; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_38 = 7'h26 == io_wa ? io_di : mem_38; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_39 = 7'h27 == io_wa ? io_di : mem_39; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_40 = 7'h28 == io_wa ? io_di : mem_40; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_41 = 7'h29 == io_wa ? io_di : mem_41; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_42 = 7'h2a == io_wa ? io_di : mem_42; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_43 = 7'h2b == io_wa ? io_di : mem_43; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_44 = 7'h2c == io_wa ? io_di : mem_44; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_45 = 7'h2d == io_wa ? io_di : mem_45; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_46 = 7'h2e == io_wa ? io_di : mem_46; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_47 = 7'h2f == io_wa ? io_di : mem_47; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_48 = 7'h30 == io_wa ? io_di : mem_48; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_49 = 7'h31 == io_wa ? io_di : mem_49; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_50 = 7'h32 == io_wa ? io_di : mem_50; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_51 = 7'h33 == io_wa ? io_di : mem_51; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_52 = 7'h34 == io_wa ? io_di : mem_52; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_53 = 7'h35 == io_wa ? io_di : mem_53; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_54 = 7'h36 == io_wa ? io_di : mem_54; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_55 = 7'h37 == io_wa ? io_di : mem_55; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_56 = 7'h38 == io_wa ? io_di : mem_56; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_57 = 7'h39 == io_wa ? io_di : mem_57; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_58 = 7'h3a == io_wa ? io_di : mem_58; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_59 = 7'h3b == io_wa ? io_di : mem_59; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_60 = 7'h3c == io_wa ? io_di : mem_60; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_61 = 7'h3d == io_wa ? io_di : mem_61; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_62 = 7'h3e == io_wa ? io_di : mem_62; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_63 = 7'h3f == io_wa ? io_di : mem_63; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_64 = 7'h40 == io_wa ? io_di : mem_64; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_65 = 7'h41 == io_wa ? io_di : mem_65; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_66 = 7'h42 == io_wa ? io_di : mem_66; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_67 = 7'h43 == io_wa ? io_di : mem_67; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_68 = 7'h44 == io_wa ? io_di : mem_68; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_69 = 7'h45 == io_wa ? io_di : mem_69; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_70 = 7'h46 == io_wa ? io_di : mem_70; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_71 = 7'h47 == io_wa ? io_di : mem_71; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_72 = 7'h48 == io_wa ? io_di : mem_72; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_73 = 7'h49 == io_wa ? io_di : mem_73; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_74 = 7'h4a == io_wa ? io_di : mem_74; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_75 = 7'h4b == io_wa ? io_di : mem_75; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_76 = 7'h4c == io_wa ? io_di : mem_76; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_77 = 7'h4d == io_wa ? io_di : mem_77; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_78 = 7'h4e == io_wa ? io_di : mem_78; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_79 = 7'h4f == io_wa ? io_di : mem_79; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_80 = 7'h50 == io_wa ? io_di : mem_80; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_81 = 7'h51 == io_wa ? io_di : mem_81; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_82 = 7'h52 == io_wa ? io_di : mem_82; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_83 = 7'h53 == io_wa ? io_di : mem_83; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_84 = 7'h54 == io_wa ? io_di : mem_84; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_85 = 7'h55 == io_wa ? io_di : mem_85; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_86 = 7'h56 == io_wa ? io_di : mem_86; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_87 = 7'h57 == io_wa ? io_di : mem_87; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_88 = 7'h58 == io_wa ? io_di : mem_88; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_89 = 7'h59 == io_wa ? io_di : mem_89; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_90 = 7'h5a == io_wa ? io_di : mem_90; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_91 = 7'h5b == io_wa ? io_di : mem_91; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_92 = 7'h5c == io_wa ? io_di : mem_92; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_93 = 7'h5d == io_wa ? io_di : mem_93; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_94 = 7'h5e == io_wa ? io_di : mem_94; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_95 = 7'h5f == io_wa ? io_di : mem_95; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_96 = 7'h60 == io_wa ? io_di : mem_96; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_97 = 7'h61 == io_wa ? io_di : mem_97; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_98 = 7'h62 == io_wa ? io_di : mem_98; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_99 = 7'h63 == io_wa ? io_di : mem_99; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_100 = 7'h64 == io_wa ? io_di : mem_100; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_101 = 7'h65 == io_wa ? io_di : mem_101; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_102 = 7'h66 == io_wa ? io_di : mem_102; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_103 = 7'h67 == io_wa ? io_di : mem_103; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_104 = 7'h68 == io_wa ? io_di : mem_104; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_105 = 7'h69 == io_wa ? io_di : mem_105; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_106 = 7'h6a == io_wa ? io_di : mem_106; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_107 = 7'h6b == io_wa ? io_di : mem_107; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_108 = 7'h6c == io_wa ? io_di : mem_108; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_109 = 7'h6d == io_wa ? io_di : mem_109; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_110 = 7'h6e == io_wa ? io_di : mem_110; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_111 = 7'h6f == io_wa ? io_di : mem_111; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_112 = 7'h70 == io_wa ? io_di : mem_112; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_113 = 7'h71 == io_wa ? io_di : mem_113; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_114 = 7'h72 == io_wa ? io_di : mem_114; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_115 = 7'h73 == io_wa ? io_di : mem_115; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_116 = 7'h74 == io_wa ? io_di : mem_116; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_117 = 7'h75 == io_wa ? io_di : mem_117; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_118 = 7'h76 == io_wa ? io_di : mem_118; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_119 = 7'h77 == io_wa ? io_di : mem_119; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_120 = 7'h78 == io_wa ? io_di : mem_120; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_121 = 7'h79 == io_wa ? io_di : mem_121; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_122 = 7'h7a == io_wa ? io_di : mem_122; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_123 = 7'h7b == io_wa ? io_di : mem_123; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_124 = 7'h7c == io_wa ? io_di : mem_124; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_125 = 7'h7d == io_wa ? io_di : mem_125; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_126 = 7'h7e == io_wa ? io_di : mem_126; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_127 = 7'h7f == io_wa ? io_di : mem_127; // @[nv_ram_rwsp.scala 37:20:@12.6]
  assign _GEN_258 = 7'h1 == ra_d ? mem_1 : mem_0; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_259 = 7'h2 == ra_d ? mem_2 : _GEN_258; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_260 = 7'h3 == ra_d ? mem_3 : _GEN_259; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_261 = 7'h4 == ra_d ? mem_4 : _GEN_260; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_262 = 7'h5 == ra_d ? mem_5 : _GEN_261; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_263 = 7'h6 == ra_d ? mem_6 : _GEN_262; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_264 = 7'h7 == ra_d ? mem_7 : _GEN_263; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_265 = 7'h8 == ra_d ? mem_8 : _GEN_264; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_266 = 7'h9 == ra_d ? mem_9 : _GEN_265; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_267 = 7'ha == ra_d ? mem_10 : _GEN_266; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_268 = 7'hb == ra_d ? mem_11 : _GEN_267; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_269 = 7'hc == ra_d ? mem_12 : _GEN_268; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_270 = 7'hd == ra_d ? mem_13 : _GEN_269; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_271 = 7'he == ra_d ? mem_14 : _GEN_270; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_272 = 7'hf == ra_d ? mem_15 : _GEN_271; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_273 = 7'h10 == ra_d ? mem_16 : _GEN_272; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_274 = 7'h11 == ra_d ? mem_17 : _GEN_273; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_275 = 7'h12 == ra_d ? mem_18 : _GEN_274; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_276 = 7'h13 == ra_d ? mem_19 : _GEN_275; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_277 = 7'h14 == ra_d ? mem_20 : _GEN_276; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_278 = 7'h15 == ra_d ? mem_21 : _GEN_277; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_279 = 7'h16 == ra_d ? mem_22 : _GEN_278; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_280 = 7'h17 == ra_d ? mem_23 : _GEN_279; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_281 = 7'h18 == ra_d ? mem_24 : _GEN_280; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_282 = 7'h19 == ra_d ? mem_25 : _GEN_281; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_283 = 7'h1a == ra_d ? mem_26 : _GEN_282; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_284 = 7'h1b == ra_d ? mem_27 : _GEN_283; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_285 = 7'h1c == ra_d ? mem_28 : _GEN_284; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_286 = 7'h1d == ra_d ? mem_29 : _GEN_285; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_287 = 7'h1e == ra_d ? mem_30 : _GEN_286; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_288 = 7'h1f == ra_d ? mem_31 : _GEN_287; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_289 = 7'h20 == ra_d ? mem_32 : _GEN_288; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_290 = 7'h21 == ra_d ? mem_33 : _GEN_289; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_291 = 7'h22 == ra_d ? mem_34 : _GEN_290; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_292 = 7'h23 == ra_d ? mem_35 : _GEN_291; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_293 = 7'h24 == ra_d ? mem_36 : _GEN_292; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_294 = 7'h25 == ra_d ? mem_37 : _GEN_293; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_295 = 7'h26 == ra_d ? mem_38 : _GEN_294; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_296 = 7'h27 == ra_d ? mem_39 : _GEN_295; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_297 = 7'h28 == ra_d ? mem_40 : _GEN_296; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_298 = 7'h29 == ra_d ? mem_41 : _GEN_297; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_299 = 7'h2a == ra_d ? mem_42 : _GEN_298; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_300 = 7'h2b == ra_d ? mem_43 : _GEN_299; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_301 = 7'h2c == ra_d ? mem_44 : _GEN_300; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_302 = 7'h2d == ra_d ? mem_45 : _GEN_301; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_303 = 7'h2e == ra_d ? mem_46 : _GEN_302; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_304 = 7'h2f == ra_d ? mem_47 : _GEN_303; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_305 = 7'h30 == ra_d ? mem_48 : _GEN_304; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_306 = 7'h31 == ra_d ? mem_49 : _GEN_305; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_307 = 7'h32 == ra_d ? mem_50 : _GEN_306; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_308 = 7'h33 == ra_d ? mem_51 : _GEN_307; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_309 = 7'h34 == ra_d ? mem_52 : _GEN_308; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_310 = 7'h35 == ra_d ? mem_53 : _GEN_309; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_311 = 7'h36 == ra_d ? mem_54 : _GEN_310; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_312 = 7'h37 == ra_d ? mem_55 : _GEN_311; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_313 = 7'h38 == ra_d ? mem_56 : _GEN_312; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_314 = 7'h39 == ra_d ? mem_57 : _GEN_313; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_315 = 7'h3a == ra_d ? mem_58 : _GEN_314; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_316 = 7'h3b == ra_d ? mem_59 : _GEN_315; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_317 = 7'h3c == ra_d ? mem_60 : _GEN_316; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_318 = 7'h3d == ra_d ? mem_61 : _GEN_317; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_319 = 7'h3e == ra_d ? mem_62 : _GEN_318; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_320 = 7'h3f == ra_d ? mem_63 : _GEN_319; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_321 = 7'h40 == ra_d ? mem_64 : _GEN_320; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_322 = 7'h41 == ra_d ? mem_65 : _GEN_321; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_323 = 7'h42 == ra_d ? mem_66 : _GEN_322; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_324 = 7'h43 == ra_d ? mem_67 : _GEN_323; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_325 = 7'h44 == ra_d ? mem_68 : _GEN_324; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_326 = 7'h45 == ra_d ? mem_69 : _GEN_325; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_327 = 7'h46 == ra_d ? mem_70 : _GEN_326; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_328 = 7'h47 == ra_d ? mem_71 : _GEN_327; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_329 = 7'h48 == ra_d ? mem_72 : _GEN_328; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_330 = 7'h49 == ra_d ? mem_73 : _GEN_329; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_331 = 7'h4a == ra_d ? mem_74 : _GEN_330; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_332 = 7'h4b == ra_d ? mem_75 : _GEN_331; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_333 = 7'h4c == ra_d ? mem_76 : _GEN_332; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_334 = 7'h4d == ra_d ? mem_77 : _GEN_333; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_335 = 7'h4e == ra_d ? mem_78 : _GEN_334; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_336 = 7'h4f == ra_d ? mem_79 : _GEN_335; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_337 = 7'h50 == ra_d ? mem_80 : _GEN_336; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_338 = 7'h51 == ra_d ? mem_81 : _GEN_337; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_339 = 7'h52 == ra_d ? mem_82 : _GEN_338; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_340 = 7'h53 == ra_d ? mem_83 : _GEN_339; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_341 = 7'h54 == ra_d ? mem_84 : _GEN_340; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_342 = 7'h55 == ra_d ? mem_85 : _GEN_341; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_343 = 7'h56 == ra_d ? mem_86 : _GEN_342; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_344 = 7'h57 == ra_d ? mem_87 : _GEN_343; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_345 = 7'h58 == ra_d ? mem_88 : _GEN_344; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_346 = 7'h59 == ra_d ? mem_89 : _GEN_345; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_347 = 7'h5a == ra_d ? mem_90 : _GEN_346; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_348 = 7'h5b == ra_d ? mem_91 : _GEN_347; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_349 = 7'h5c == ra_d ? mem_92 : _GEN_348; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_350 = 7'h5d == ra_d ? mem_93 : _GEN_349; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_351 = 7'h5e == ra_d ? mem_94 : _GEN_350; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_352 = 7'h5f == ra_d ? mem_95 : _GEN_351; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_353 = 7'h60 == ra_d ? mem_96 : _GEN_352; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_354 = 7'h61 == ra_d ? mem_97 : _GEN_353; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_355 = 7'h62 == ra_d ? mem_98 : _GEN_354; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_356 = 7'h63 == ra_d ? mem_99 : _GEN_355; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_357 = 7'h64 == ra_d ? mem_100 : _GEN_356; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_358 = 7'h65 == ra_d ? mem_101 : _GEN_357; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_359 = 7'h66 == ra_d ? mem_102 : _GEN_358; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_360 = 7'h67 == ra_d ? mem_103 : _GEN_359; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_361 = 7'h68 == ra_d ? mem_104 : _GEN_360; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_362 = 7'h69 == ra_d ? mem_105 : _GEN_361; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_363 = 7'h6a == ra_d ? mem_106 : _GEN_362; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_364 = 7'h6b == ra_d ? mem_107 : _GEN_363; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_365 = 7'h6c == ra_d ? mem_108 : _GEN_364; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_366 = 7'h6d == ra_d ? mem_109 : _GEN_365; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_367 = 7'h6e == ra_d ? mem_110 : _GEN_366; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_368 = 7'h6f == ra_d ? mem_111 : _GEN_367; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_369 = 7'h70 == ra_d ? mem_112 : _GEN_368; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_370 = 7'h71 == ra_d ? mem_113 : _GEN_369; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_371 = 7'h72 == ra_d ? mem_114 : _GEN_370; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_372 = 7'h73 == ra_d ? mem_115 : _GEN_371; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_373 = 7'h74 == ra_d ? mem_116 : _GEN_372; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_374 = 7'h75 == ra_d ? mem_117 : _GEN_373; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_375 = 7'h76 == ra_d ? mem_118 : _GEN_374; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_376 = 7'h77 == ra_d ? mem_119 : _GEN_375; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_377 = 7'h78 == ra_d ? mem_120 : _GEN_376; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_378 = 7'h79 == ra_d ? mem_121 : _GEN_377; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_379 = 7'h7a == ra_d ? mem_122 : _GEN_378; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_380 = 7'h7b == ra_d ? mem_123 : _GEN_379; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_381 = 7'h7c == ra_d ? mem_124 : _GEN_380; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_382 = 7'h7d == ra_d ? mem_125 : _GEN_381; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_383 = 7'h7e == ra_d ? mem_126 : _GEN_382; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign _GEN_384 = 7'h7f == ra_d ? mem_127 : _GEN_383; // @[nv_ram_rwsp.scala 44:16:@18.6]
  assign io_dout = dout_r; // @[nv_ram_rwsp.scala 46:13:@20.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mem_0 = _RAND_0[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_1 = _RAND_1[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_2 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mem_3 = _RAND_3[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_4 = _RAND_4[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_5 = _RAND_5[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mem_6 = _RAND_6[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_7 = _RAND_7[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_8 = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mem_9 = _RAND_9[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_10 = _RAND_10[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_11 = _RAND_11[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mem_12 = _RAND_12[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mem_13 = _RAND_13[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mem_14 = _RAND_14[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mem_15 = _RAND_15[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mem_16 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mem_17 = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mem_18 = _RAND_18[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mem_19 = _RAND_19[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mem_20 = _RAND_20[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  mem_21 = _RAND_21[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_22 = _RAND_22[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_23 = _RAND_23[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_24 = _RAND_24[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_25 = _RAND_25[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_26 = _RAND_26[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_27 = _RAND_27[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_28 = _RAND_28[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_29 = _RAND_29[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_30 = _RAND_30[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_31 = _RAND_31[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_32 = _RAND_32[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  mem_33 = _RAND_33[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  mem_34 = _RAND_34[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  mem_35 = _RAND_35[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mem_36 = _RAND_36[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  mem_37 = _RAND_37[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mem_38 = _RAND_38[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  mem_39 = _RAND_39[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  mem_40 = _RAND_40[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  mem_41 = _RAND_41[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  mem_42 = _RAND_42[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  mem_43 = _RAND_43[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  mem_44 = _RAND_44[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  mem_45 = _RAND_45[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  mem_46 = _RAND_46[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  mem_47 = _RAND_47[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  mem_48 = _RAND_48[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  mem_49 = _RAND_49[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  mem_50 = _RAND_50[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  mem_51 = _RAND_51[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  mem_52 = _RAND_52[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  mem_53 = _RAND_53[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  mem_54 = _RAND_54[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  mem_55 = _RAND_55[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  mem_56 = _RAND_56[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  mem_57 = _RAND_57[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  mem_58 = _RAND_58[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  mem_59 = _RAND_59[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  mem_60 = _RAND_60[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  mem_61 = _RAND_61[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  mem_62 = _RAND_62[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  mem_63 = _RAND_63[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  mem_64 = _RAND_64[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  mem_65 = _RAND_65[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_66 = _RAND_66[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  mem_67 = _RAND_67[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  mem_68 = _RAND_68[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  mem_69 = _RAND_69[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  mem_70 = _RAND_70[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  mem_71 = _RAND_71[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  mem_72 = _RAND_72[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  mem_73 = _RAND_73[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  mem_74 = _RAND_74[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  mem_75 = _RAND_75[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  mem_76 = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  mem_77 = _RAND_77[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  mem_78 = _RAND_78[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  mem_79 = _RAND_79[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  mem_80 = _RAND_80[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  mem_81 = _RAND_81[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  mem_82 = _RAND_82[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  mem_83 = _RAND_83[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  mem_84 = _RAND_84[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  mem_85 = _RAND_85[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  mem_86 = _RAND_86[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  mem_87 = _RAND_87[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  mem_88 = _RAND_88[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  mem_89 = _RAND_89[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  mem_90 = _RAND_90[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  mem_91 = _RAND_91[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  mem_92 = _RAND_92[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  mem_93 = _RAND_93[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  mem_94 = _RAND_94[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  mem_95 = _RAND_95[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  mem_96 = _RAND_96[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  mem_97 = _RAND_97[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  mem_98 = _RAND_98[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  mem_99 = _RAND_99[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  mem_100 = _RAND_100[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  mem_101 = _RAND_101[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  mem_102 = _RAND_102[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  mem_103 = _RAND_103[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  mem_104 = _RAND_104[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  mem_105 = _RAND_105[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  mem_106 = _RAND_106[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  mem_107 = _RAND_107[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  mem_108 = _RAND_108[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  mem_109 = _RAND_109[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  mem_110 = _RAND_110[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  mem_111 = _RAND_111[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  mem_112 = _RAND_112[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  mem_113 = _RAND_113[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  mem_114 = _RAND_114[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  mem_115 = _RAND_115[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  mem_116 = _RAND_116[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  mem_117 = _RAND_117[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  mem_118 = _RAND_118[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  mem_119 = _RAND_119[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  mem_120 = _RAND_120[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  mem_121 = _RAND_121[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  mem_122 = _RAND_122[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  mem_123 = _RAND_123[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  mem_124 = _RAND_124[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  mem_125 = _RAND_125[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  mem_126 = _RAND_126[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  mem_127 = _RAND_127[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  ra_d = _RAND_128[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  dout_r = _RAND_129[10:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_clk) begin
    if (io_we) begin
      if (7'h0 == io_wa) begin
        mem_0 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1 == io_wa) begin
        mem_1 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2 == io_wa) begin
        mem_2 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3 == io_wa) begin
        mem_3 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4 == io_wa) begin
        mem_4 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5 == io_wa) begin
        mem_5 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6 == io_wa) begin
        mem_6 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7 == io_wa) begin
        mem_7 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h8 == io_wa) begin
        mem_8 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h9 == io_wa) begin
        mem_9 <= io_di;
      end
    end
    if (io_we) begin
      if (7'ha == io_wa) begin
        mem_10 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hb == io_wa) begin
        mem_11 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hc == io_wa) begin
        mem_12 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hd == io_wa) begin
        mem_13 <= io_di;
      end
    end
    if (io_we) begin
      if (7'he == io_wa) begin
        mem_14 <= io_di;
      end
    end
    if (io_we) begin
      if (7'hf == io_wa) begin
        mem_15 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h10 == io_wa) begin
        mem_16 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h11 == io_wa) begin
        mem_17 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h12 == io_wa) begin
        mem_18 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h13 == io_wa) begin
        mem_19 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h14 == io_wa) begin
        mem_20 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h15 == io_wa) begin
        mem_21 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h16 == io_wa) begin
        mem_22 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h17 == io_wa) begin
        mem_23 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h18 == io_wa) begin
        mem_24 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h19 == io_wa) begin
        mem_25 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1a == io_wa) begin
        mem_26 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1b == io_wa) begin
        mem_27 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1c == io_wa) begin
        mem_28 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1d == io_wa) begin
        mem_29 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1e == io_wa) begin
        mem_30 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h1f == io_wa) begin
        mem_31 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h20 == io_wa) begin
        mem_32 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h21 == io_wa) begin
        mem_33 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h22 == io_wa) begin
        mem_34 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h23 == io_wa) begin
        mem_35 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h24 == io_wa) begin
        mem_36 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h25 == io_wa) begin
        mem_37 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h26 == io_wa) begin
        mem_38 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h27 == io_wa) begin
        mem_39 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h28 == io_wa) begin
        mem_40 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h29 == io_wa) begin
        mem_41 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2a == io_wa) begin
        mem_42 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2b == io_wa) begin
        mem_43 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2c == io_wa) begin
        mem_44 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2d == io_wa) begin
        mem_45 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2e == io_wa) begin
        mem_46 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h2f == io_wa) begin
        mem_47 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h30 == io_wa) begin
        mem_48 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h31 == io_wa) begin
        mem_49 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h32 == io_wa) begin
        mem_50 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h33 == io_wa) begin
        mem_51 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h34 == io_wa) begin
        mem_52 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h35 == io_wa) begin
        mem_53 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h36 == io_wa) begin
        mem_54 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h37 == io_wa) begin
        mem_55 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h38 == io_wa) begin
        mem_56 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h39 == io_wa) begin
        mem_57 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3a == io_wa) begin
        mem_58 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3b == io_wa) begin
        mem_59 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3c == io_wa) begin
        mem_60 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3d == io_wa) begin
        mem_61 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3e == io_wa) begin
        mem_62 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h3f == io_wa) begin
        mem_63 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h40 == io_wa) begin
        mem_64 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h41 == io_wa) begin
        mem_65 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h42 == io_wa) begin
        mem_66 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h43 == io_wa) begin
        mem_67 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h44 == io_wa) begin
        mem_68 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h45 == io_wa) begin
        mem_69 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h46 == io_wa) begin
        mem_70 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h47 == io_wa) begin
        mem_71 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h48 == io_wa) begin
        mem_72 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h49 == io_wa) begin
        mem_73 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4a == io_wa) begin
        mem_74 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4b == io_wa) begin
        mem_75 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4c == io_wa) begin
        mem_76 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4d == io_wa) begin
        mem_77 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4e == io_wa) begin
        mem_78 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h4f == io_wa) begin
        mem_79 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h50 == io_wa) begin
        mem_80 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h51 == io_wa) begin
        mem_81 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h52 == io_wa) begin
        mem_82 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h53 == io_wa) begin
        mem_83 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h54 == io_wa) begin
        mem_84 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h55 == io_wa) begin
        mem_85 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h56 == io_wa) begin
        mem_86 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h57 == io_wa) begin
        mem_87 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h58 == io_wa) begin
        mem_88 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h59 == io_wa) begin
        mem_89 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5a == io_wa) begin
        mem_90 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5b == io_wa) begin
        mem_91 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5c == io_wa) begin
        mem_92 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5d == io_wa) begin
        mem_93 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5e == io_wa) begin
        mem_94 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h5f == io_wa) begin
        mem_95 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h60 == io_wa) begin
        mem_96 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h61 == io_wa) begin
        mem_97 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h62 == io_wa) begin
        mem_98 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h63 == io_wa) begin
        mem_99 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h64 == io_wa) begin
        mem_100 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h65 == io_wa) begin
        mem_101 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h66 == io_wa) begin
        mem_102 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h67 == io_wa) begin
        mem_103 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h68 == io_wa) begin
        mem_104 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h69 == io_wa) begin
        mem_105 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6a == io_wa) begin
        mem_106 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6b == io_wa) begin
        mem_107 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6c == io_wa) begin
        mem_108 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6d == io_wa) begin
        mem_109 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6e == io_wa) begin
        mem_110 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h6f == io_wa) begin
        mem_111 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h70 == io_wa) begin
        mem_112 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h71 == io_wa) begin
        mem_113 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h72 == io_wa) begin
        mem_114 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h73 == io_wa) begin
        mem_115 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h74 == io_wa) begin
        mem_116 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h75 == io_wa) begin
        mem_117 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h76 == io_wa) begin
        mem_118 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h77 == io_wa) begin
        mem_119 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h78 == io_wa) begin
        mem_120 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h79 == io_wa) begin
        mem_121 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7a == io_wa) begin
        mem_122 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7b == io_wa) begin
        mem_123 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7c == io_wa) begin
        mem_124 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7d == io_wa) begin
        mem_125 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7e == io_wa) begin
        mem_126 <= io_di;
      end
    end
    if (io_we) begin
      if (7'h7f == io_wa) begin
        mem_127 <= io_di;
      end
    end
    if (io_re) begin
      ra_d <= io_ra;
    end
    if (io_ore) begin
      if (7'h7f == ra_d) begin
        dout_r <= mem_127;
      end else begin
        if (7'h7e == ra_d) begin
          dout_r <= mem_126;
        end else begin
          if (7'h7d == ra_d) begin
            dout_r <= mem_125;
          end else begin
            if (7'h7c == ra_d) begin
              dout_r <= mem_124;
            end else begin
              if (7'h7b == ra_d) begin
                dout_r <= mem_123;
              end else begin
                if (7'h7a == ra_d) begin
                  dout_r <= mem_122;
                end else begin
                  if (7'h79 == ra_d) begin
                    dout_r <= mem_121;
                  end else begin
                    if (7'h78 == ra_d) begin
                      dout_r <= mem_120;
                    end else begin
                      if (7'h77 == ra_d) begin
                        dout_r <= mem_119;
                      end else begin
                        if (7'h76 == ra_d) begin
                          dout_r <= mem_118;
                        end else begin
                          if (7'h75 == ra_d) begin
                            dout_r <= mem_117;
                          end else begin
                            if (7'h74 == ra_d) begin
                              dout_r <= mem_116;
                            end else begin
                              if (7'h73 == ra_d) begin
                                dout_r <= mem_115;
                              end else begin
                                if (7'h72 == ra_d) begin
                                  dout_r <= mem_114;
                                end else begin
                                  if (7'h71 == ra_d) begin
                                    dout_r <= mem_113;
                                  end else begin
                                    if (7'h70 == ra_d) begin
                                      dout_r <= mem_112;
                                    end else begin
                                      if (7'h6f == ra_d) begin
                                        dout_r <= mem_111;
                                      end else begin
                                        if (7'h6e == ra_d) begin
                                          dout_r <= mem_110;
                                        end else begin
                                          if (7'h6d == ra_d) begin
                                            dout_r <= mem_109;
                                          end else begin
                                            if (7'h6c == ra_d) begin
                                              dout_r <= mem_108;
                                            end else begin
                                              if (7'h6b == ra_d) begin
                                                dout_r <= mem_107;
                                              end else begin
                                                if (7'h6a == ra_d) begin
                                                  dout_r <= mem_106;
                                                end else begin
                                                  if (7'h69 == ra_d) begin
                                                    dout_r <= mem_105;
                                                  end else begin
                                                    if (7'h68 == ra_d) begin
                                                      dout_r <= mem_104;
                                                    end else begin
                                                      if (7'h67 == ra_d) begin
                                                        dout_r <= mem_103;
                                                      end else begin
                                                        if (7'h66 == ra_d) begin
                                                          dout_r <= mem_102;
                                                        end else begin
                                                          if (7'h65 == ra_d) begin
                                                            dout_r <= mem_101;
                                                          end else begin
                                                            if (7'h64 == ra_d) begin
                                                              dout_r <= mem_100;
                                                            end else begin
                                                              if (7'h63 == ra_d) begin
                                                                dout_r <= mem_99;
                                                              end else begin
                                                                if (7'h62 == ra_d) begin
                                                                  dout_r <= mem_98;
                                                                end else begin
                                                                  if (7'h61 == ra_d) begin
                                                                    dout_r <= mem_97;
                                                                  end else begin
                                                                    if (7'h60 == ra_d) begin
                                                                      dout_r <= mem_96;
                                                                    end else begin
                                                                      if (7'h5f == ra_d) begin
                                                                        dout_r <= mem_95;
                                                                      end else begin
                                                                        if (7'h5e == ra_d) begin
                                                                          dout_r <= mem_94;
                                                                        end else begin
                                                                          if (7'h5d == ra_d) begin
                                                                            dout_r <= mem_93;
                                                                          end else begin
                                                                            if (7'h5c == ra_d) begin
                                                                              dout_r <= mem_92;
                                                                            end else begin
                                                                              if (7'h5b == ra_d) begin
                                                                                dout_r <= mem_91;
                                                                              end else begin
                                                                                if (7'h5a == ra_d) begin
                                                                                  dout_r <= mem_90;
                                                                                end else begin
                                                                                  if (7'h59 == ra_d) begin
                                                                                    dout_r <= mem_89;
                                                                                  end else begin
                                                                                    if (7'h58 == ra_d) begin
                                                                                      dout_r <= mem_88;
                                                                                    end else begin
                                                                                      if (7'h57 == ra_d) begin
                                                                                        dout_r <= mem_87;
                                                                                      end else begin
                                                                                        if (7'h56 == ra_d) begin
                                                                                          dout_r <= mem_86;
                                                                                        end else begin
                                                                                          if (7'h55 == ra_d) begin
                                                                                            dout_r <= mem_85;
                                                                                          end else begin
                                                                                            if (7'h54 == ra_d) begin
                                                                                              dout_r <= mem_84;
                                                                                            end else begin
                                                                                              if (7'h53 == ra_d) begin
                                                                                                dout_r <= mem_83;
                                                                                              end else begin
                                                                                                if (7'h52 == ra_d) begin
                                                                                                  dout_r <= mem_82;
                                                                                                end else begin
                                                                                                  if (7'h51 == ra_d) begin
                                                                                                    dout_r <= mem_81;
                                                                                                  end else begin
                                                                                                    if (7'h50 == ra_d) begin
                                                                                                      dout_r <= mem_80;
                                                                                                    end else begin
                                                                                                      if (7'h4f == ra_d) begin
                                                                                                        dout_r <= mem_79;
                                                                                                      end else begin
                                                                                                        if (7'h4e == ra_d) begin
                                                                                                          dout_r <= mem_78;
                                                                                                        end else begin
                                                                                                          if (7'h4d == ra_d) begin
                                                                                                            dout_r <= mem_77;
                                                                                                          end else begin
                                                                                                            if (7'h4c == ra_d) begin
                                                                                                              dout_r <= mem_76;
                                                                                                            end else begin
                                                                                                              if (7'h4b == ra_d) begin
                                                                                                                dout_r <= mem_75;
                                                                                                              end else begin
                                                                                                                if (7'h4a == ra_d) begin
                                                                                                                  dout_r <= mem_74;
                                                                                                                end else begin
                                                                                                                  if (7'h49 == ra_d) begin
                                                                                                                    dout_r <= mem_73;
                                                                                                                  end else begin
                                                                                                                    if (7'h48 == ra_d) begin
                                                                                                                      dout_r <= mem_72;
                                                                                                                    end else begin
                                                                                                                      if (7'h47 == ra_d) begin
                                                                                                                        dout_r <= mem_71;
                                                                                                                      end else begin
                                                                                                                        if (7'h46 == ra_d) begin
                                                                                                                          dout_r <= mem_70;
                                                                                                                        end else begin
                                                                                                                          if (7'h45 == ra_d) begin
                                                                                                                            dout_r <= mem_69;
                                                                                                                          end else begin
                                                                                                                            if (7'h44 == ra_d) begin
                                                                                                                              dout_r <= mem_68;
                                                                                                                            end else begin
                                                                                                                              if (7'h43 == ra_d) begin
                                                                                                                                dout_r <= mem_67;
                                                                                                                              end else begin
                                                                                                                                if (7'h42 == ra_d) begin
                                                                                                                                  dout_r <= mem_66;
                                                                                                                                end else begin
                                                                                                                                  if (7'h41 == ra_d) begin
                                                                                                                                    dout_r <= mem_65;
                                                                                                                                  end else begin
                                                                                                                                    if (7'h40 == ra_d) begin
                                                                                                                                      dout_r <= mem_64;
                                                                                                                                    end else begin
                                                                                                                                      if (7'h3f == ra_d) begin
                                                                                                                                        dout_r <= mem_63;
                                                                                                                                      end else begin
                                                                                                                                        if (7'h3e == ra_d) begin
                                                                                                                                          dout_r <= mem_62;
                                                                                                                                        end else begin
                                                                                                                                          if (7'h3d == ra_d) begin
                                                                                                                                            dout_r <= mem_61;
                                                                                                                                          end else begin
                                                                                                                                            if (7'h3c == ra_d) begin
                                                                                                                                              dout_r <= mem_60;
                                                                                                                                            end else begin
                                                                                                                                              if (7'h3b == ra_d) begin
                                                                                                                                                dout_r <= mem_59;
                                                                                                                                              end else begin
                                                                                                                                                if (7'h3a == ra_d) begin
                                                                                                                                                  dout_r <= mem_58;
                                                                                                                                                end else begin
                                                                                                                                                  if (7'h39 == ra_d) begin
                                                                                                                                                    dout_r <= mem_57;
                                                                                                                                                  end else begin
                                                                                                                                                    if (7'h38 == ra_d) begin
                                                                                                                                                      dout_r <= mem_56;
                                                                                                                                                    end else begin
                                                                                                                                                      if (7'h37 == ra_d) begin
                                                                                                                                                        dout_r <= mem_55;
                                                                                                                                                      end else begin
                                                                                                                                                        if (7'h36 == ra_d) begin
                                                                                                                                                          dout_r <= mem_54;
                                                                                                                                                        end else begin
                                                                                                                                                          if (7'h35 == ra_d) begin
                                                                                                                                                            dout_r <= mem_53;
                                                                                                                                                          end else begin
                                                                                                                                                            if (7'h34 == ra_d) begin
                                                                                                                                                              dout_r <= mem_52;
                                                                                                                                                            end else begin
                                                                                                                                                              if (7'h33 == ra_d) begin
                                                                                                                                                                dout_r <= mem_51;
                                                                                                                                                              end else begin
                                                                                                                                                                if (7'h32 == ra_d) begin
                                                                                                                                                                  dout_r <= mem_50;
                                                                                                                                                                end else begin
                                                                                                                                                                  if (7'h31 == ra_d) begin
                                                                                                                                                                    dout_r <= mem_49;
                                                                                                                                                                  end else begin
                                                                                                                                                                    if (7'h30 == ra_d) begin
                                                                                                                                                                      dout_r <= mem_48;
                                                                                                                                                                    end else begin
                                                                                                                                                                      if (7'h2f == ra_d) begin
                                                                                                                                                                        dout_r <= mem_47;
                                                                                                                                                                      end else begin
                                                                                                                                                                        if (7'h2e == ra_d) begin
                                                                                                                                                                          dout_r <= mem_46;
                                                                                                                                                                        end else begin
                                                                                                                                                                          if (7'h2d == ra_d) begin
                                                                                                                                                                            dout_r <= mem_45;
                                                                                                                                                                          end else begin
                                                                                                                                                                            if (7'h2c == ra_d) begin
                                                                                                                                                                              dout_r <= mem_44;
                                                                                                                                                                            end else begin
                                                                                                                                                                              if (7'h2b == ra_d) begin
                                                                                                                                                                                dout_r <= mem_43;
                                                                                                                                                                              end else begin
                                                                                                                                                                                if (7'h2a == ra_d) begin
                                                                                                                                                                                  dout_r <= mem_42;
                                                                                                                                                                                end else begin
                                                                                                                                                                                  if (7'h29 == ra_d) begin
                                                                                                                                                                                    dout_r <= mem_41;
                                                                                                                                                                                  end else begin
                                                                                                                                                                                    if (7'h28 == ra_d) begin
                                                                                                                                                                                      dout_r <= mem_40;
                                                                                                                                                                                    end else begin
                                                                                                                                                                                      if (7'h27 == ra_d) begin
                                                                                                                                                                                        dout_r <= mem_39;
                                                                                                                                                                                      end else begin
                                                                                                                                                                                        if (7'h26 == ra_d) begin
                                                                                                                                                                                          dout_r <= mem_38;
                                                                                                                                                                                        end else begin
                                                                                                                                                                                          if (7'h25 == ra_d) begin
                                                                                                                                                                                            dout_r <= mem_37;
                                                                                                                                                                                          end else begin
                                                                                                                                                                                            if (7'h24 == ra_d) begin
                                                                                                                                                                                              dout_r <= mem_36;
                                                                                                                                                                                            end else begin
                                                                                                                                                                                              if (7'h23 == ra_d) begin
                                                                                                                                                                                                dout_r <= mem_35;
                                                                                                                                                                                              end else begin
                                                                                                                                                                                                if (7'h22 == ra_d) begin
                                                                                                                                                                                                  dout_r <= mem_34;
                                                                                                                                                                                                end else begin
                                                                                                                                                                                                  if (7'h21 == ra_d) begin
                                                                                                                                                                                                    dout_r <= mem_33;
                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                    if (7'h20 == ra_d) begin
                                                                                                                                                                                                      dout_r <= mem_32;
                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                      if (7'h1f == ra_d) begin
                                                                                                                                                                                                        dout_r <= mem_31;
                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                        if (7'h1e == ra_d) begin
                                                                                                                                                                                                          dout_r <= mem_30;
                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                          if (7'h1d == ra_d) begin
                                                                                                                                                                                                            dout_r <= mem_29;
                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                            if (7'h1c == ra_d) begin
                                                                                                                                                                                                              dout_r <= mem_28;
                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                              if (7'h1b == ra_d) begin
                                                                                                                                                                                                                dout_r <= mem_27;
                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                if (7'h1a == ra_d) begin
                                                                                                                                                                                                                  dout_r <= mem_26;
                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                  if (7'h19 == ra_d) begin
                                                                                                                                                                                                                    dout_r <= mem_25;
                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                    if (7'h18 == ra_d) begin
                                                                                                                                                                                                                      dout_r <= mem_24;
                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                      if (7'h17 == ra_d) begin
                                                                                                                                                                                                                        dout_r <= mem_23;
                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                        if (7'h16 == ra_d) begin
                                                                                                                                                                                                                          dout_r <= mem_22;
                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                          if (7'h15 == ra_d) begin
                                                                                                                                                                                                                            dout_r <= mem_21;
                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                            if (7'h14 == ra_d) begin
                                                                                                                                                                                                                              dout_r <= mem_20;
                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                              if (7'h13 == ra_d) begin
                                                                                                                                                                                                                                dout_r <= mem_19;
                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                if (7'h12 == ra_d) begin
                                                                                                                                                                                                                                  dout_r <= mem_18;
                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                  if (7'h11 == ra_d) begin
                                                                                                                                                                                                                                    dout_r <= mem_17;
                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                    if (7'h10 == ra_d) begin
                                                                                                                                                                                                                                      dout_r <= mem_16;
                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                      if (7'hf == ra_d) begin
                                                                                                                                                                                                                                        dout_r <= mem_15;
                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                        if (7'he == ra_d) begin
                                                                                                                                                                                                                                          dout_r <= mem_14;
                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                          if (7'hd == ra_d) begin
                                                                                                                                                                                                                                            dout_r <= mem_13;
                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                            if (7'hc == ra_d) begin
                                                                                                                                                                                                                                              dout_r <= mem_12;
                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                              if (7'hb == ra_d) begin
                                                                                                                                                                                                                                                dout_r <= mem_11;
                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                if (7'ha == ra_d) begin
                                                                                                                                                                                                                                                  dout_r <= mem_10;
                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                  if (7'h9 == ra_d) begin
                                                                                                                                                                                                                                                    dout_r <= mem_9;
                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                    if (7'h8 == ra_d) begin
                                                                                                                                                                                                                                                      dout_r <= mem_8;
                                                                                                                                                                                                                                                    end else begin
                                                                                                                                                                                                                                                      if (7'h7 == ra_d) begin
                                                                                                                                                                                                                                                        dout_r <= mem_7;
                                                                                                                                                                                                                                                      end else begin
                                                                                                                                                                                                                                                        if (7'h6 == ra_d) begin
                                                                                                                                                                                                                                                          dout_r <= mem_6;
                                                                                                                                                                                                                                                        end else begin
                                                                                                                                                                                                                                                          if (7'h5 == ra_d) begin
                                                                                                                                                                                                                                                            dout_r <= mem_5;
                                                                                                                                                                                                                                                          end else begin
                                                                                                                                                                                                                                                            if (7'h4 == ra_d) begin
                                                                                                                                                                                                                                                              dout_r <= mem_4;
                                                                                                                                                                                                                                                            end else begin
                                                                                                                                                                                                                                                              if (7'h3 == ra_d) begin
                                                                                                                                                                                                                                                                dout_r <= mem_3;
                                                                                                                                                                                                                                                              end else begin
                                                                                                                                                                                                                                                                if (7'h2 == ra_d) begin
                                                                                                                                                                                                                                                                  dout_r <= mem_2;
                                                                                                                                                                                                                                                                end else begin
                                                                                                                                                                                                                                                                  if (7'h1 == ra_d) begin
                                                                                                                                                                                                                                                                    dout_r <= mem_1;
                                                                                                                                                                                                                                                                  end else begin
                                                                                                                                                                                                                                                                    dout_r <= mem_0;
                                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                                end
                                                                                                                                                                                                                                              end
                                                                                                                                                                                                                                            end
                                                                                                                                                                                                                                          end
                                                                                                                                                                                                                                        end
                                                                                                                                                                                                                                      end
                                                                                                                                                                                                                                    end
                                                                                                                                                                                                                                  end
                                                                                                                                                                                                                                end
                                                                                                                                                                                                                              end
                                                                                                                                                                                                                            end
                                                                                                                                                                                                                          end
                                                                                                                                                                                                                        end
                                                                                                                                                                                                                      end
                                                                                                                                                                                                                    end
                                                                                                                                                                                                                  end
                                                                                                                                                                                                                end
                                                                                                                                                                                                              end
                                                                                                                                                                                                            end
                                                                                                                                                                                                          end
                                                                                                                                                                                                        end
                                                                                                                                                                                                      end
                                                                                                                                                                                                    end
                                                                                                                                                                                                  end
                                                                                                                                                                                                end
                                                                                                                                                                                              end
                                                                                                                                                                                            end
                                                                                                                                                                                          end
                                                                                                                                                                                        end
                                                                                                                                                                                      end
                                                                                                                                                                                    end
                                                                                                                                                                                  end
                                                                                                                                                                                end
                                                                                                                                                                              end
                                                                                                                                                                            end
                                                                                                                                                                          end
                                                                                                                                                                        end
                                                                                                                                                                      end
                                                                                                                                                                    end
                                                                                                                                                                  end
                                                                                                                                                                end
                                                                                                                                                              end
                                                                                                                                                            end
                                                                                                                                                          end
                                                                                                                                                        end
                                                                                                                                                      end
                                                                                                                                                    end
                                                                                                                                                  end
                                                                                                                                                end
                                                                                                                                              end
                                                                                                                                            end
                                                                                                                                          end
                                                                                                                                        end
                                                                                                                                      end
                                                                                                                                    end
                                                                                                                                  end
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
  end
endmodule

module NV_soDLA_CSC_dl_for_check( // @[:@3.2]
  input          nvdla_core_clk, // @[:@6.4]
  input          nvdla_core_ng_clk, // @[:@6.4]
  input          nvdla_core_rstn, // @[:@6.4]
  input  [1:0]   sc_state, // @[:@6.4]
  input          sg2dl_reuse_rls, // @[:@6.4]
  input          sg2dl_pvld, // @[:@6.4]
  input  [30:0]  sg2dl_pd, // @[:@6.4]
  input          cdma2sc_dat_updt, // @[:@6.4]
  input  [14:0]  cdma2sc_dat_entries, // @[:@6.4]
  input  [13:0]  cdma2sc_dat_slices, // @[:@6.4]
  input          sc2cdma_dat_pending_req, // @[:@6.4]
  output         sc2cdma_dat_updt, // @[:@6.4]
  output [14:0]  sc2cdma_dat_entries, // @[:@6.4]
  output [13:0]  sc2cdma_dat_slices, // @[:@6.4]

  output         sc2buf_dat_rd_en, // @[:@6.4]
  output [12:0]  sc2buf_dat_rd_addr, // @[:@6.4]

  input          sc2buf_dat_rd_valid, // @[:@6.4]
  input  [511:0] sc2buf_dat_rd_data, // @[:@6.4]


  output         sc2mac_dat_a_valid, // @[:@6.4]
  output [63:0]  sc2mac_dat_a_mask, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data0, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data1, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data2, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data3, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data4, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data5, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data6, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data7, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data8, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data9, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data10, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data11, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data12, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data13, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data14, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data15, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data16, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data17, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data18, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data19, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data20, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data21, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data22, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data23, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data24, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data25, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data26, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data27, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data28, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data29, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data30, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data31, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data32, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data33, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data34, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data35, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data36, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data37, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data38, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data39, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data40, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data41, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data42, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data43, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data44, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data45, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data46, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data47, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data48, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data49, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data50, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data51, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data52, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data53, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data54, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data55, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data56, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data57, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data58, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data59, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data60, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data61, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data62, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data63, // @[:@6.4]
  output [8:0]   sc2mac_dat_a_pd, // @[:@6.4]
  output         sc2mac_dat_b_valid, // @[:@6.4]
  output [63:0]  sc2mac_dat_b_mask, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data0, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data1, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data2, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data3, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data4, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data5, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data6, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data7, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data8, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data9, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data10, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data11, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data12, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data13, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data14, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data15, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data16, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data17, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data18, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data19, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data20, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data21, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data22, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data23, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data24, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data25, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data26, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data27, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data28, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data29, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data30, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data31, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data32, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data33, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data34, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data35, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data36, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data37, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data38, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data39, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data40, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data41, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data42, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data43, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data44, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data45, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data46, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data47, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data48, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data49, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data50, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data51, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data52, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data53, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data54, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data55, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data56, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data57, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data58, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data59, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data60, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data61, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data62, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data63, // @[:@6.4]
  output [8:0]   sc2mac_dat_b_pd, // @[:@6.4]
  input          reg2dp_op_en, // @[:@6.4]
  input          reg2dp_conv_mode, // @[:@6.4]
  input  [4:0]   reg2dp_batches, // @[:@6.4]
  input  [1:0]   reg2dp_proc_precision, // @[:@6.4]
  input          reg2dp_datain_format, // @[:@6.4]
  input          reg2dp_skip_data_rls, // @[:@6.4]
  input  [12:0]  reg2dp_datain_channel_ext, // @[:@6.4]
  input  [12:0]  reg2dp_datain_height_ext, // @[:@6.4]
  input  [12:0]  reg2dp_datain_width_ext, // @[:@6.4]
  input  [1:0]   reg2dp_y_extension, // @[:@6.4]
  input  [12:0]  reg2dp_weight_channel_ext, // @[:@6.4]
  input  [13:0]  reg2dp_entries, // @[:@6.4]
  input  [12:0]  reg2dp_dataout_width, // @[:@6.4]
  input  [11:0]  reg2dp_rls_slices, // @[:@6.4]
  input  [2:0]   reg2dp_conv_x_stride_ext, // @[:@6.4]
  input  [2:0]   reg2dp_conv_y_stride_ext, // @[:@6.4]
  input  [4:0]   reg2dp_x_dilation_ext, // @[:@6.4]
  input  [4:0]   reg2dp_y_dilation_ext, // @[:@6.4]
  input  [4:0]   reg2dp_pad_left, // @[:@6.4]
  input  [4:0]   reg2dp_pad_top, // @[:@6.4]
  input  [15:0]  reg2dp_pad_value, // @[:@6.4]
  input  [4:0]   reg2dp_data_bank, // @[:@6.4]
  input  [1:0]   reg2dp_pra_truncate, // @[:@6.4]
  output         slcg_wg_en // @[:@6.4]
);
  wire  _T_337; // @[NV_NVDLA_CSC_dl_for_check.scala 95:38:@8.4]
  wire  _T_339; // @[NV_NVDLA_CSC_dl_for_check.scala 99:31:@9.4]
  wire  _T_343; // @[NV_NVDLA_CSC_dl_for_check.scala 101:31:@11.4]
  wire  _T_347; // @[NV_NVDLA_CSC_dl_for_check.scala 108:32:@14.4]
  wire  _T_351; // @[NV_NVDLA_CSC_dl_for_check.scala 110:35:@16.4]
  wire  _T_352; // @[NV_NVDLA_CSC_dl_for_check.scala 111:22:@17.4]
  wire [6:0] _T_357; // @[NV_NVDLA_CSC_dl_for_check.scala 118:53:@18.4]
  wire [6:0] _T_359; // @[NV_NVDLA_CSC_dl_for_check.scala 118:24:@19.4]
  wire [2:0] _T_360; // @[NV_NVDLA_CSC_dl_for_check.scala 118:100:@20.4]
  wire [2:0] _T_362; // @[NV_NVDLA_CSC_dl_for_check.scala 119:22:@21.4]
  wire [3:0] _T_364; // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@22.4]
  wire [3:0] _T_365; // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@23.4]
  wire [3:0] _T_367; // @[NV_NVDLA_CSC_dl_for_check.scala 121:51:@24.4]
  wire [1:0] _T_368; // @[NV_NVDLA_CSC_dl_for_check.scala 122:62:@25.4]
  wire [5:0] _T_371; // @[Cat.scala 30:58:@26.4]
  wire [4:0] _T_374; // @[Cat.scala 30:58:@27.4]
  wire [4:0] _GEN_671; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  wire [5:0] _T_375; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  wire  _T_376; // @[Mux.scala 46:19:@29.4]
  wire [5:0] _T_377; // @[Mux.scala 46:16:@30.4]
  wire  _T_378; // @[Mux.scala 46:19:@31.4]
  wire [5:0] _T_379; // @[Mux.scala 46:16:@32.4]
  wire  _T_381; // @[NV_NVDLA_CSC_dl_for_check.scala 126:88:@33.4]
  wire [5:0] _T_387; // @[NV_NVDLA_CSC_dl_for_check.scala 126:172:@35.4]
  wire [5:0] _T_388; // @[NV_NVDLA_CSC_dl_for_check.scala 126:58:@36.4]
  wire [6:0] _T_391; // @[Cat.scala 30:58:@37.4]
  wire [6:0] _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  wire [7:0] _T_392; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  wire [6:0] _T_393; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@39.4]
  wire [6:0] _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  wire [7:0] _T_395; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  wire [6:0] _T_396; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@42.4]
  wire [6:0] _T_399; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@44.4]
  wire [5:0] _T_400; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@45.4]
  wire  _T_401; // @[Mux.scala 46:19:@46.4]
  wire [5:0] _T_402; // @[Mux.scala 46:16:@47.4]
  wire  _T_403; // @[Mux.scala 46:19:@48.4]
  wire [6:0] _T_404; // @[Mux.scala 46:16:@49.4]
  wire [6:0] _T_407; // @[NV_NVDLA_CSC_dl_for_check.scala 129:80:@51.4]
  wire [7:0] _T_410; // @[Cat.scala 30:58:@52.4]
  wire [6:0] _T_415; // @[Mux.scala 46:16:@55.4]
  wire [7:0] _T_417; // @[Mux.scala 46:16:@57.4]
  wire [11:0] _T_419; // @[Cat.scala 30:58:@58.4]
  wire [3:0] _T_421; // @[NV_NVDLA_CSC_dl_for_check.scala 139:52:@59.4]
  wire [5:0] _T_424; // @[NV_NVDLA_CSC_dl_for_check.scala 140:60:@60.4]
  wire [5:0] _T_425; // @[NV_NVDLA_CSC_dl_for_check.scala 140:21:@61.4]
  wire [5:0] _T_428; // @[NV_NVDLA_CSC_dl_for_check.scala 141:60:@62.4]
  wire [5:0] _T_429; // @[NV_NVDLA_CSC_dl_for_check.scala 141:21:@63.4]
  reg  _T_432; // @[NV_NVDLA_CSC_dl_for_check.scala 143:26:@64.4]
  reg [31:0] _RAND_0;
  reg [5:0] _T_439; // @[NV_NVDLA_CSC_dl_for_check.scala 144:25:@66.4]
  reg [31:0] _RAND_1;
  reg [13:0] _T_446; // @[NV_NVDLA_CSC_dl_for_check.scala 145:25:@68.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_453; // @[NV_NVDLA_CSC_dl_for_check.scala 146:29:@70.4]
  reg [31:0] _RAND_3;
  reg [14:0] _T_460; // @[NV_NVDLA_CSC_dl_for_check.scala 147:22:@72.4]
  reg [31:0] _RAND_4;
  reg [14:0] _T_467; // @[NV_NVDLA_CSC_dl_for_check.scala 148:28:@74.4]
  reg [31:0] _RAND_5;
  reg [12:0] _T_474; // @[NV_NVDLA_CSC_dl_for_check.scala 149:32:@76.4]
  reg [31:0] _RAND_6;
  reg [14:0] _T_488; // @[NV_NVDLA_CSC_dl_for_check.scala 151:26:@80.4]
  reg [31:0] _RAND_7;
  reg [11:0] _T_495; // @[NV_NVDLA_CSC_dl_for_check.scala 152:30:@82.4]
  reg [31:0] _RAND_8;
  reg [11:0] _T_502; // @[NV_NVDLA_CSC_dl_for_check.scala 153:30:@84.4]
  reg [31:0] _RAND_9;
  reg [13:0] _T_509; // @[NV_NVDLA_CSC_dl_for_check.scala 154:25:@86.4]
  reg [31:0] _RAND_10;
  wire [14:0] _T_511; // @[NV_NVDLA_CSC_dl_for_check.scala 157:43:@87.4]
  wire [20:0] _T_513; // @[NV_NVDLA_CSC_dl_for_check.scala 158:41:@89.4]
  wire [14:0] _T_514; // @[NV_NVDLA_CSC_dl_for_check.scala 158:56:@90.4]
  wire [11:0] _T_515; // @[NV_NVDLA_CSC_dl_for_check.scala 160:37:@91.4]
  wire [14:0] _GEN_674; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  wire [20:0] _T_516; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  wire [11:0] _T_517; // @[NV_NVDLA_CSC_dl_for_check.scala 161:47:@93.4]
  wire [14:0] _GEN_675; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  wire [28:0] _T_518; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  wire [11:0] _T_519; // @[NV_NVDLA_CSC_dl_for_check.scala 162:51:@95.4]
  wire [12:0] _T_521; // @[NV_NVDLA_CSC_dl_for_check.scala 163:41:@96.4]
  wire [11:0] _T_522; // @[NV_NVDLA_CSC_dl_for_check.scala 163:41:@97.4]
  wire [13:0] _T_524; // @[NV_NVDLA_CSC_dl_for_check.scala 164:77:@98.4]
  wire [12:0] _GEN_676; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@99.4]
  wire [13:0] _T_525; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@99.4]
  wire [13:0] _T_526; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@100.4]
  wire [13:0] _T_527; // @[NV_NVDLA_CSC_dl_for_check.scala 164:23:@101.4]
  wire [13:0] _T_528; // @[NV_NVDLA_CSC_dl_for_check.scala 165:24:@102.4]
  wire [14:0] _GEN_677; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@103.4]
  wire [28:0] _T_529; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@103.4]
  wire [14:0] _T_530; // @[NV_NVDLA_CSC_dl_for_check.scala 166:54:@104.4]
  reg [33:0] _T_548; // @[NV_NVDLA_CSC_dl_for_check.scala 171:24:@110.4]
  reg [63:0] _RAND_11;
  reg [4:0] _T_555; // @[NV_NVDLA_CSC_dl_for_check.scala 172:24:@112.4]
  reg [31:0] _RAND_12;
  reg [13:0] _T_562; // @[NV_NVDLA_CSC_dl_for_check.scala 173:27:@114.4]
  reg [31:0] _RAND_13;
  reg [12:0] _T_569; // @[NV_NVDLA_CSC_dl_for_check.scala 174:31:@116.4]
  reg [31:0] _RAND_14;
  reg [12:0] _T_576; // @[NV_NVDLA_CSC_dl_for_check.scala 175:32:@118.4]
  reg [31:0] _RAND_15;
  reg [10:0] _T_583; // @[NV_NVDLA_CSC_dl_for_check.scala 176:33:@120.4]
  reg [31:0] _RAND_16;
  reg [2:0] _T_586; // @[NV_NVDLA_CSC_dl_for_check.scala 177:29:@121.4]
  reg [31:0] _RAND_17;
  reg [2:0] _T_589; // @[NV_NVDLA_CSC_dl_for_check.scala 178:29:@122.4]
  reg [31:0] _RAND_18;
  reg [2:0] _T_595; // @[NV_NVDLA_CSC_dl_for_check.scala 180:29:@124.4]
  reg [31:0] _RAND_19;
  reg [2:0] _T_598; // @[NV_NVDLA_CSC_dl_for_check.scala 181:29:@125.4]
  reg [31:0] _RAND_20;
  reg [2:0] _T_601; // @[NV_NVDLA_CSC_dl_for_check.scala 182:29:@126.4]
  reg [31:0] _RAND_21;
  reg [2:0] _T_604; // @[NV_NVDLA_CSC_dl_for_check.scala 183:29:@127.4]
  reg [31:0] _RAND_22;
  reg [2:0] _T_610; // @[NV_NVDLA_CSC_dl_for_check.scala 185:29:@129.4]
  reg [31:0] _RAND_23;
  reg [2:0] _T_613; // @[NV_NVDLA_CSC_dl_for_check.scala 186:29:@130.4]
  reg [31:0] _RAND_24;
  reg [2:0] _T_619; // @[NV_NVDLA_CSC_dl_for_check.scala 188:30:@132.4]
  reg [31:0] _RAND_25;
  reg [2:0] _T_622; // @[NV_NVDLA_CSC_dl_for_check.scala 189:27:@133.4]
  reg [31:0] _RAND_26;
  reg [2:0] _T_625; // @[NV_NVDLA_CSC_dl_for_check.scala 190:27:@134.4]
  reg [31:0] _RAND_27;
  reg [3:0] _T_632; // @[NV_NVDLA_CSC_dl_for_check.scala 191:28:@136.4]
  reg [31:0] _RAND_28;
  reg [3:0] _T_639; // @[NV_NVDLA_CSC_dl_for_check.scala 192:28:@138.4]
  reg [31:0] _RAND_29;
  reg [4:0] _T_649; // @[NV_NVDLA_CSC_dl_for_check.scala 194:24:@141.4]
  reg [31:0] _RAND_30;
  reg [6:0] _T_656; // @[NV_NVDLA_CSC_dl_for_check.scala 195:27:@143.4]
  reg [31:0] _RAND_31;
  reg [6:0] _T_663; // @[NV_NVDLA_CSC_dl_for_check.scala 196:34:@145.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_670; // @[NV_NVDLA_CSC_dl_for_check.scala 197:26:@147.4]
  reg [31:0] _RAND_33;
  reg [6:0] _T_677; // @[NV_NVDLA_CSC_dl_for_check.scala 198:34:@149.4]
  reg [31:0] _RAND_34;
  reg [11:0] _T_684; // @[NV_NVDLA_CSC_dl_for_check.scala 199:30:@151.4]
  reg [31:0] _RAND_35;
  reg [5:0] _T_691; // @[NV_NVDLA_CSC_dl_for_check.scala 200:23:@153.4]
  reg [31:0] _RAND_36;
  reg [5:0] _T_698; // @[NV_NVDLA_CSC_dl_for_check.scala 201:23:@155.4]
  reg [31:0] _RAND_37;
  reg [15:0] _T_705; // @[NV_NVDLA_CSC_dl_for_check.scala 202:24:@157.4]
  reg [31:0] _RAND_38;
  reg [14:0] _T_712; // @[NV_NVDLA_CSC_dl_for_check.scala 203:26:@159.4]
  reg [31:0] _RAND_39;
  reg [14:0] _T_719; // @[NV_NVDLA_CSC_dl_for_check.scala 204:30:@161.4]
  reg [31:0] _RAND_40;
  reg [14:0] _T_726; // @[NV_NVDLA_CSC_dl_for_check.scala 205:30:@163.4]
  reg [31:0] _RAND_41;
  reg [13:0] _T_733; // @[NV_NVDLA_CSC_dl_for_check.scala 207:26:@165.4]
  reg [31:0] _RAND_42;
  reg [14:0] _T_740; // @[NV_NVDLA_CSC_dl_for_check.scala 208:27:@167.4]
  reg [31:0] _RAND_43;
  wire [33:0] _T_755; // @[Bitwise.scala 72:12:@175.6]
  wire [5:0] _T_757; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@177.6]
  wire [4:0] _T_758; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@178.6]
  wire [13:0] _T_760; // @[NV_NVDLA_CSC_dl_for_check.scala 216:48:@180.6]
  wire [6:0] _T_766; // @[NV_NVDLA_CSC_dl_for_check.scala 219:93:@185.6]
  wire [10:0] _T_767; // @[Cat.scala 30:58:@186.6]
  wire [14:0] _T_771; // @[Cat.scala 30:58:@219.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [4:0] _GEN_2; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [13:0] _GEN_3; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [12:0] _GEN_4; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [12:0] _GEN_5; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [10:0] _GEN_6; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_7; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_8; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_10; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_11; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_12; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_13; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_15; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_19; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [2:0] _GEN_20; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [3:0] _GEN_21; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [5:0] _GEN_24; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [6:0] _GEN_26; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [6:0] _GEN_27; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [11:0] _GEN_30; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [5:0] _GEN_31; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [14:0] _GEN_34; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [14:0] _GEN_35; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [14:0] _GEN_36; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [13:0] _GEN_37; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [13:0] _GEN_39; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [12:0] _GEN_40; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  wire [11:0] _GEN_43; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  wire [11:0] _GEN_44; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  wire [14:0] _GEN_45; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  wire [14:0] _GEN_46; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  wire [14:0] _GEN_47; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  wire [13:0] _GEN_48; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@239.4]
  wire [14:0] _GEN_49; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@239.4]
  reg [14:0] _T_793; // @[NV_NVDLA_CSC_dl_for_check.scala 287:59:@251.4]
  reg [31:0] _RAND_44;
  wire  _T_873; // @[NV_NVDLA_CSC_dl_for_check.scala 328:37:@314.4]
  wire  _T_874; // @[NV_NVDLA_CSC_dl_for_check.scala 328:23:@315.4]
  wire  _T_1958; // @[NV_NVDLA_CSC_dl_for_check.scala 918:32:@1229.4]
  reg  _T_1934; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1197.4]
  reg [31:0] _RAND_45;
  wire  _T_1959; // @[NV_NVDLA_CSC_dl_for_check.scala 918:36:@1230.4]
  wire  _T_1960; // @[NV_NVDLA_CSC_dl_for_check.scala 919:35:@1231.4]
  reg  _T_1928; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1195.4]
  reg [31:0] _RAND_46;
  wire  _T_1961; // @[NV_NVDLA_CSC_dl_for_check.scala 919:39:@1232.4]
  wire  _T_1962; // @[NV_NVDLA_CSC_dl_for_check.scala 918:57:@1233.4]
  wire  _T_1963; // @[NV_NVDLA_CSC_dl_for_check.scala 920:35:@1234.4]
  reg  _T_1925; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1194.4]
  reg [31:0] _RAND_47;
  wire  _T_1964; // @[NV_NVDLA_CSC_dl_for_check.scala 920:39:@1235.4]
  wire  _T_1965; // @[NV_NVDLA_CSC_dl_for_check.scala 919:60:@1236.4]
  wire  _T_1966; // @[NV_NVDLA_CSC_dl_for_check.scala 927:42:@1238.4]
  wire [26:0] _T_1970; // @[Bitwise.scala 72:12:@1240.4]
  reg [26:0] _T_1948; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1202.4]
  reg [31:0] _RAND_48;
  wire [26:0] _T_1971; // @[NV_NVDLA_CSC_dl_for_check.scala 927:47:@1241.4]
  wire  _T_1972; // @[NV_NVDLA_CSC_dl_for_check.scala 928:42:@1242.4]
  wire [26:0] _T_1976; // @[Bitwise.scala 72:12:@1244.4]
  reg [26:0] _T_1942; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1200.4]
  reg [31:0] _RAND_49;
  wire [26:0] _T_1977; // @[NV_NVDLA_CSC_dl_for_check.scala 928:47:@1245.4]
  wire [26:0] _T_1978; // @[NV_NVDLA_CSC_dl_for_check.scala 927:66:@1246.4]
  wire  _T_1979; // @[NV_NVDLA_CSC_dl_for_check.scala 929:42:@1247.4]
  wire [26:0] _T_1983; // @[Bitwise.scala 72:12:@1249.4]
  reg [26:0] _T_1939; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1199.4]
  reg [31:0] _RAND_50;
  wire [26:0] _T_1984; // @[NV_NVDLA_CSC_dl_for_check.scala 929:47:@1250.4]
  wire [26:0] _T_1985; // @[NV_NVDLA_CSC_dl_for_check.scala 928:66:@1251.4]
  wire  _T_2004; // @[NV_NVDLA_CSC_dl_for_check.scala 953:26:@1270.4]
  wire  _T_871; // @[NV_NVDLA_CSC_dl_for_check.scala 325:29:@313.4]
  wire  _T_876; // @[NV_NVDLA_CSC_dl_for_check.scala 328:66:@316.4]
  wire  _T_877; // @[NV_NVDLA_CSC_dl_for_check.scala 328:53:@317.4]
  wire  _T_878; // @[NV_NVDLA_CSC_dl_for_check.scala 328:42:@318.4]
  wire [13:0] _T_879; // @[NV_NVDLA_CSC_dl_for_check.scala 329:28:@320.4]
  wire [14:0] _T_880; // @[NV_NVDLA_CSC_dl_for_check.scala 330:29:@322.4]
  wire [14:0] _T_811; // @[NV_NVDLA_CSC_dl_for_check.scala 297:28:@262.4]
  wire [15:0] _T_819; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@269.4]
  wire [14:0] _T_820; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@270.4]
  wire [13:0] _T_826; // @[Cat.scala 30:58:@272.4]
  wire [14:0] _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@273.4]
  wire [15:0] _T_827; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@273.4]
  wire [15:0] _T_828; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@274.4]
  wire [14:0] _T_829; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@275.4]
  wire  _T_836; // @[NV_NVDLA_CSC_dl_for_check.scala 304:45:@278.4]
  wire [14:0] _T_838; // @[NV_NVDLA_CSC_dl_for_check.scala 305:83:@279.4]
  wire [14:0] _T_839; // @[NV_NVDLA_CSC_dl_for_check.scala 305:25:@280.4]
  wire  _T_865; // @[NV_NVDLA_CSC_dl_for_check.scala 316:13:@303.4]
  wire [14:0] _GEN_52; // @[NV_NVDLA_CSC_dl_for_check.scala 316:25:@304.4]
  reg  _T_883; // @[NV_NVDLA_CSC_dl_for_check.scala 332:31:@324.4]
  reg [31:0] _RAND_51;
  reg [13:0] _T_886; // @[Reg.scala 19:20:@327.4]
  reg [31:0] _RAND_52;
  wire [13:0] _GEN_54; // @[Reg.scala 20:19:@328.4]
  reg [14:0] _T_889; // @[Reg.scala 19:20:@332.4]
  reg [31:0] _RAND_53;
  wire [14:0] _GEN_55; // @[Reg.scala 20:19:@333.4]
  reg  _T_894; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@338.4]
  reg [31:0] _RAND_54;
  reg  _T_897; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@339.4]
  reg [31:0] _RAND_55;
  reg  _T_900; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@340.4]
  reg [31:0] _RAND_56;
  reg  _T_903; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@341.4]
  reg [31:0] _RAND_57;
  reg  _T_906; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@342.4]
  reg [31:0] _RAND_58;
  reg  _T_928; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@372.4]
  reg [31:0] _RAND_59;
  reg  _T_931; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@373.4]
  reg [31:0] _RAND_60;
  reg  _T_934; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@374.4]
  reg [31:0] _RAND_61;
  reg  _T_937; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@375.4]
  reg [31:0] _RAND_62;
  reg [30:0] _T_942; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@377.4]
  reg [31:0] _RAND_63;
  reg [30:0] _T_945; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@378.4]
  reg [31:0] _RAND_64;
  reg [30:0] _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@379.4]
  reg [31:0] _RAND_65;
  reg [30:0] _T_951; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@380.4]
  reg [31:0] _RAND_66;
  wire [30:0] _T_939; // @[NV_NVDLA_CSC_dl_for_check.scala 365:19:@376.4 NV_NVDLA_CSC_dl_for_check.scala 369:12:@382.4]
  wire [30:0] _GEN_61; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@384.4]
  wire [30:0] _GEN_62; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@388.4]
  wire [30:0] _GEN_63; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@392.4]
  wire [30:0] _GEN_64; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@396.4]
  wire  _T_952; // @[NV_NVDLA_CSC_dl_for_check.scala 378:30:@399.4]
  wire  _T_953; // @[NV_NVDLA_CSC_dl_for_check.scala 378:34:@400.4]
  wire  _T_954; // @[NV_NVDLA_CSC_dl_for_check.scala 379:30:@401.4]
  wire  _T_955; // @[NV_NVDLA_CSC_dl_for_check.scala 379:34:@402.4]
  wire  _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 378:50:@403.4]
  wire  _T_957; // @[NV_NVDLA_CSC_dl_for_check.scala 380:30:@404.4]
  wire  _T_958; // @[NV_NVDLA_CSC_dl_for_check.scala 380:34:@405.4]
  wire  _T_959; // @[NV_NVDLA_CSC_dl_for_check.scala 379:50:@406.4]
  wire  _T_960; // @[NV_NVDLA_CSC_dl_for_check.scala 382:37:@407.4]
  wire [30:0] _T_964; // @[Bitwise.scala 72:12:@409.4]
  wire [30:0] _T_965; // @[NV_NVDLA_CSC_dl_for_check.scala 382:42:@410.4]
  wire  _T_966; // @[NV_NVDLA_CSC_dl_for_check.scala 383:37:@411.4]
  wire [30:0] _T_970; // @[Bitwise.scala 72:12:@413.4]
  wire [30:0] _T_971; // @[NV_NVDLA_CSC_dl_for_check.scala 383:42:@414.4]
  wire [30:0] _T_972; // @[NV_NVDLA_CSC_dl_for_check.scala 382:56:@415.4]
  wire  _T_973; // @[NV_NVDLA_CSC_dl_for_check.scala 384:37:@416.4]
  wire [30:0] _T_977; // @[Bitwise.scala 72:12:@418.4]
  wire [30:0] _T_978; // @[NV_NVDLA_CSC_dl_for_check.scala 384:42:@419.4]
  wire [30:0] _T_979; // @[NV_NVDLA_CSC_dl_for_check.scala 383:56:@420.4]
  wire [4:0] _T_980; // @[NV_NVDLA_CSC_dl_for_check.scala 387:24:@421.4]
  wire [4:0] _T_981; // @[NV_NVDLA_CSC_dl_for_check.scala 388:24:@422.4]
  wire [6:0] _T_982; // @[NV_NVDLA_CSC_dl_for_check.scala 389:28:@423.4]
  wire [6:0] _T_983; // @[NV_NVDLA_CSC_dl_for_check.scala 390:29:@424.4]
  wire [1:0] _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 391:25:@425.4]
  wire  _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 392:25:@426.4]
  wire  _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 393:27:@427.4]
  wire  _T_987; // @[NV_NVDLA_CSC_dl_for_check.scala 394:25:@428.4]
  wire  _T_988; // @[NV_NVDLA_CSC_dl_for_check.scala 395:25:@429.4]
  wire  _T_989; // @[NV_NVDLA_CSC_dl_for_check.scala 396:27:@430.4]
  reg [4:0] _T_996; // @[NV_NVDLA_CSC_dl_for_check.scala 401:24:@433.4]
  reg [31:0] _RAND_67;
  wire [5:0] _T_1000; // @[NV_NVDLA_CSC_dl_for_check.scala 405:24:@434.4]
  wire [4:0] _T_1001; // @[NV_NVDLA_CSC_dl_for_check.scala 405:24:@435.4]
  wire  _T_1004; // @[NV_NVDLA_CSC_dl_for_check.scala 407:27:@439.4]
  wire [4:0] _T_1002; // @[NV_NVDLA_CSC_dl_for_check.scala 404:17:@436.4]
  wire [4:0] _T_1003; // @[NV_NVDLA_CSC_dl_for_check.scala 403:17:@437.4]
  reg [1:0] _T_1007; // @[NV_NVDLA_CSC_dl_for_check.scala 410:24:@441.4]
  reg [31:0] _RAND_68;
  wire [2:0] _T_1011; // @[NV_NVDLA_CSC_dl_for_check.scala 413:31:@443.4]
  wire [1:0] _T_1012; // @[NV_NVDLA_CSC_dl_for_check.scala 413:31:@444.4]
  wire [2:0] _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 414:32:@445.4]
  wire  _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 414:32:@445.4]
  wire  _T_1015; // @[NV_NVDLA_CSC_dl_for_check.scala 415:61:@447.4]
  reg [6:0] _T_1023; // @[NV_NVDLA_CSC_dl_for_check.scala 421:25:@455.4]
  reg [31:0] _RAND_69;
  wire  _T_1063; // @[NV_NVDLA_CSC_dl_for_check.scala 448:37:@484.4]
  wire  _T_1064; // @[NV_NVDLA_CSC_dl_for_check.scala 448:24:@485.4]
  wire  _T_1066; // @[NV_NVDLA_CSC_dl_for_check.scala 448:56:@486.4]
  wire  _T_1067; // @[NV_NVDLA_CSC_dl_for_check.scala 448:44:@487.4]
  wire  _T_1068; // @[NV_NVDLA_CSC_dl_for_check.scala 448:42:@488.4]
  wire  _T_1070; // @[NV_NVDLA_CSC_dl_for_check.scala 448:75:@489.4]
  wire  _T_1071; // @[NV_NVDLA_CSC_dl_for_check.scala 448:63:@490.4]
  wire  _T_1072; // @[NV_NVDLA_CSC_dl_for_check.scala 448:61:@491.4]
  reg  _T_1052; // @[NV_NVDLA_CSC_dl_for_check.scala 440:32:@477.4]
  reg [31:0] _RAND_70;
  wire  _T_1074; // @[NV_NVDLA_CSC_dl_for_check.scala 448:22:@492.4]
  wire  _T_1075; // @[NV_NVDLA_CSC_dl_for_check.scala 447:22:@493.4]
  wire  _T_1016; // @[NV_NVDLA_CSC_dl_for_check.scala 415:66:@448.4]
  wire  _T_1017; // @[NV_NVDLA_CSC_dl_for_check.scala 415:33:@449.4]
  wire  _T_1018; // @[NV_NVDLA_CSC_dl_for_check.scala 417:31:@451.6]
  wire [1:0] _T_1020; // @[NV_NVDLA_CSC_dl_for_check.scala 417:21:@452.6]
  wire [1:0] _GEN_65; // @[NV_NVDLA_CSC_dl_for_check.scala 416:23:@450.4]
  wire [7:0] _T_1029; // @[NV_NVDLA_CSC_dl_for_check.scala 425:33:@458.4]
  wire [6:0] _T_1030; // @[NV_NVDLA_CSC_dl_for_check.scala 425:33:@459.4]
  wire  _T_1031; // @[NV_NVDLA_CSC_dl_for_check.scala 426:51:@460.4]
  wire  _T_1032; // @[NV_NVDLA_CSC_dl_for_check.scala 426:33:@461.4]
  wire  _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 427:34:@463.4]
  wire  _T_1034; // @[NV_NVDLA_CSC_dl_for_check.scala 428:52:@465.4]
  wire  _T_1035; // @[NV_NVDLA_CSC_dl_for_check.scala 428:34:@466.4]
  wire  _T_1037; // @[NV_NVDLA_CSC_dl_for_check.scala 432:41:@468.6]
  wire  _T_1038; // @[NV_NVDLA_CSC_dl_for_check.scala 432:39:@469.6]
  wire [6:0] _T_1041; // @[NV_NVDLA_CSC_dl_for_check.scala 433:22:@470.6]
  wire [6:0] _T_1042; // @[NV_NVDLA_CSC_dl_for_check.scala 432:22:@471.6]
  wire [6:0] _T_1043; // @[NV_NVDLA_CSC_dl_for_check.scala 431:22:@472.6]
  wire [6:0] _GEN_66; // @[NV_NVDLA_CSC_dl_for_check.scala 430:24:@467.4]
  reg  _T_1046; // @[NV_NVDLA_CSC_dl_for_check.scala 438:35:@475.4]
  reg [31:0] _RAND_71;
  reg  _T_1049; // @[NV_NVDLA_CSC_dl_for_check.scala 439:32:@476.4]
  reg [31:0] _RAND_72;
  wire  _T_1060; // @[NV_NVDLA_CSC_dl_for_check.scala 446:27:@482.4]
  wire  _T_1055; // @[NV_NVDLA_CSC_dl_for_check.scala 443:49:@479.4]
  wire  _T_1058; // @[NV_NVDLA_CSC_dl_for_check.scala 444:32:@480.4]
  wire  _T_1059; // @[NV_NVDLA_CSC_dl_for_check.scala 443:33:@481.4]
  reg [7:0] _T_1078; // @[NV_NVDLA_CSC_dl_for_check.scala 456:31:@498.4]
  reg [31:0] _RAND_73;
  wire [7:0] _T_1080; // @[Cat.scala 30:58:@499.4]
  wire [7:0] _GEN_67; // @[NV_NVDLA_CSC_dl_for_check.scala 458:21:@500.4]
  reg [12:0] _T_1083; // @[NV_NVDLA_CSC_dl_for_check.scala 464:28:@503.4]
  reg [31:0] _RAND_74;
  reg [12:0] _T_1086; // @[NV_NVDLA_CSC_dl_for_check.scala 465:28:@504.4]
  reg [31:0] _RAND_75;
  wire [12:0] _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@505.4]
  wire [13:0] _T_1087; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@505.4]
  wire [12:0] _T_1088; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@506.4]
  wire  _T_1089; // @[NV_NVDLA_CSC_dl_for_check.scala 469:29:@507.4]
  wire  _T_1090; // @[NV_NVDLA_CSC_dl_for_check.scala 469:61:@508.4]
  wire  _T_1091; // @[NV_NVDLA_CSC_dl_for_check.scala 469:44:@509.4]
  wire  _T_1094; // @[NV_NVDLA_CSC_dl_for_check.scala 472:43:@512.4]
  wire  _T_1095; // @[NV_NVDLA_CSC_dl_for_check.scala 472:41:@513.4]
  wire [12:0] _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 473:26:@514.4]
  wire [12:0] _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 472:26:@515.4]
  wire [12:0] _T_1098; // @[NV_NVDLA_CSC_dl_for_check.scala 471:26:@516.4]
  wire  _T_1100; // @[NV_NVDLA_CSC_dl_for_check.scala 474:70:@518.4]
  wire  _T_1101; // @[NV_NVDLA_CSC_dl_for_check.scala 474:37:@519.4]
  wire  _T_1102; // @[NV_NVDLA_CSC_dl_for_check.scala 475:55:@520.4]
  wire  _T_1103; // @[NV_NVDLA_CSC_dl_for_check.scala 475:71:@521.4]
  wire  _T_1104; // @[NV_NVDLA_CSC_dl_for_check.scala 475:37:@522.4]
  wire [12:0] _GEN_68; // @[NV_NVDLA_CSC_dl_for_check.scala 477:27:@523.4]
  wire [12:0] _GEN_69; // @[NV_NVDLA_CSC_dl_for_check.scala 480:27:@526.4]
  reg [10:0] _T_1107; // @[NV_NVDLA_CSC_dl_for_check.scala 485:27:@529.4]
  reg [31:0] _RAND_76;
  wire  _T_1108; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@530.4]
  wire  _T_1110; // @[NV_NVDLA_CSC_dl_for_check.scala 488:70:@532.4]
  wire  _T_1111; // @[NV_NVDLA_CSC_dl_for_check.scala 488:36:@533.4]
  wire [11:0] _T_1115; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@535.6]
  wire [10:0] _T_1116; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@536.6]
  wire [10:0] _T_1117; // @[NV_NVDLA_CSC_dl_for_check.scala 492:24:@537.6]
  wire [10:0] _T_1118; // @[NV_NVDLA_CSC_dl_for_check.scala 491:24:@538.6]
  wire [10:0] _GEN_70; // @[NV_NVDLA_CSC_dl_for_check.scala 490:26:@534.4]
  reg [13:0] _T_1121; // @[NV_NVDLA_CSC_dl_for_check.scala 497:27:@541.4]
  reg [31:0] _RAND_77;
  reg [13:0] _T_1124; // @[NV_NVDLA_CSC_dl_for_check.scala 498:27:@542.4]
  reg [31:0] _RAND_78;
  reg [15:0] _T_1127; // @[NV_NVDLA_CSC_dl_for_check.scala 499:26:@543.4]
  reg [31:0] _RAND_79;
  reg [15:0] _T_1130; // @[NV_NVDLA_CSC_dl_for_check.scala 500:26:@544.4]
  reg [31:0] _RAND_80;
  reg [15:0] _T_1133; // @[NV_NVDLA_CSC_dl_for_check.scala 501:29:@545.4]
  reg [31:0] _RAND_81;
  reg [12:0] _T_1136; // @[NV_NVDLA_CSC_dl_for_check.scala 502:29:@546.4]
  reg [31:0] _RAND_82;
  reg  _T_1141; // @[NV_NVDLA_CSC_dl_for_check.scala 504:33:@548.4]
  reg [31:0] _RAND_83;
  reg  _T_1144; // @[NV_NVDLA_CSC_dl_for_check.scala 505:35:@549.4]
  reg [31:0] _RAND_84;
  wire [12:0] _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@550.4]
  wire [13:0] _T_1147; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@550.4]
  wire [13:0] _T_1148; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@551.4]
  wire [13:0] _T_1149; // @[NV_NVDLA_CSC_dl_for_check.scala 507:26:@552.4]
  wire [13:0] _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@553.4]
  wire [14:0] _T_1150; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@553.4]
  wire [13:0] _T_1151; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@554.4]
  wire [13:0] _T_1154; // @[NV_NVDLA_CSC_dl_for_check.scala 514:25:@557.4]
  wire [13:0] _T_1155; // @[NV_NVDLA_CSC_dl_for_check.scala 513:25:@558.4]
  wire [13:0] _T_1156; // @[NV_NVDLA_CSC_dl_for_check.scala 512:25:@559.4]
  wire [5:0] _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@560.4]
  wire [10:0] _T_1157; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@560.4]
  wire [13:0] _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 517:33:@561.4]
  wire [14:0] _T_1158; // @[NV_NVDLA_CSC_dl_for_check.scala 517:33:@561.4]
  wire [13:0] _T_1159; // @[NV_NVDLA_CSC_dl_for_check.scala 517:33:@562.4]
  wire  _T_1162; // @[NV_NVDLA_CSC_dl_for_check.scala 518:96:@565.4]
  wire  _T_1163; // @[NV_NVDLA_CSC_dl_for_check.scala 518:86:@566.4]
  wire  _T_1164; // @[NV_NVDLA_CSC_dl_for_check.scala 518:84:@567.4]
  wire  _T_1165; // @[NV_NVDLA_CSC_dl_for_check.scala 518:36:@568.4]
  wire  _T_1168; // @[NV_NVDLA_CSC_dl_for_check.scala 519:99:@571.4]
  wire  _T_1169; // @[NV_NVDLA_CSC_dl_for_check.scala 519:89:@572.4]
  wire  _T_1170; // @[NV_NVDLA_CSC_dl_for_check.scala 519:87:@573.4]
  wire  _T_1171; // @[NV_NVDLA_CSC_dl_for_check.scala 519:36:@574.4]
  wire [7:0] _T_1173; // @[NV_NVDLA_CSC_dl_for_check.scala 522:26:@575.4]
  wire  _T_1176; // @[NV_NVDLA_CSC_dl_for_check.scala 524:79:@577.4]
  wire [7:0] _T_1180; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@580.4]
  wire [6:0] _T_1181; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@581.4]
  wire [6:0] _T_1182; // @[NV_NVDLA_CSC_dl_for_check.scala 524:27:@582.4]
  wire  _T_1183; // @[NV_NVDLA_CSC_dl_for_check.scala 526:37:@583.4]
  wire  _T_1185; // @[NV_NVDLA_CSC_dl_for_check.scala 527:35:@584.4]
  wire [13:0] _T_1187; // @[NV_NVDLA_CSC_dl_for_check.scala 527:66:@585.4]
  wire [12:0] _T_1188; // @[NV_NVDLA_CSC_dl_for_check.scala 527:66:@586.4]
  wire [12:0] _T_1189; // @[NV_NVDLA_CSC_dl_for_check.scala 527:22:@587.4]
  wire [12:0] _T_1190; // @[NV_NVDLA_CSC_dl_for_check.scala 526:22:@588.4]
  wire [12:0] _GEN_688; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@590.4]
  wire  _T_1191; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@590.4]
  wire  _T_1192; // @[NV_NVDLA_CSC_dl_for_check.scala 533:39:@591.4]
  wire  _T_1193; // @[NV_NVDLA_CSC_dl_for_check.scala 533:54:@592.4]
  wire  _T_1194; // @[NV_NVDLA_CSC_dl_for_check.scala 533:71:@593.4]
  wire  _T_1197; // @[NV_NVDLA_CSC_dl_for_check.scala 534:73:@596.4]
  wire  _T_1198; // @[NV_NVDLA_CSC_dl_for_check.scala 534:71:@597.4]
  wire [15:0] _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@598.4]
  wire [16:0] _T_1199; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@598.4]
  wire [15:0] _T_1200; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@599.4]
  wire  _T_1202; // @[NV_NVDLA_CSC_dl_for_check.scala 535:54:@601.4]
  wire [15:0] _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@602.4]
  wire [16:0] _T_1203; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@602.4]
  wire [15:0] _T_1204; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@603.4]
  wire  _T_1206; // @[NV_NVDLA_CSC_dl_for_check.scala 536:56:@605.4]
  wire  _T_1207; // @[NV_NVDLA_CSC_dl_for_check.scala 536:54:@606.4]
  wire [16:0] _T_1209; // @[NV_NVDLA_CSC_dl_for_check.scala 536:91:@607.4]
  wire [15:0] _T_1210; // @[NV_NVDLA_CSC_dl_for_check.scala 536:91:@608.4]
  wire  _T_1211; // @[NV_NVDLA_CSC_dl_for_check.scala 537:41:@609.4]
  wire  _T_1212; // @[NV_NVDLA_CSC_dl_for_check.scala 537:39:@610.4]
  wire [15:0] _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@611.4]
  wire [16:0] _T_1213; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@611.4]
  wire [15:0] _T_1214; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@612.4]
  wire [15:0] _T_1215; // @[NV_NVDLA_CSC_dl_for_check.scala 537:24:@613.4]
  wire [15:0] _T_1216; // @[NV_NVDLA_CSC_dl_for_check.scala 536:24:@614.4]
  wire [15:0] _T_1217; // @[NV_NVDLA_CSC_dl_for_check.scala 535:24:@615.4]
  wire [15:0] _T_1218; // @[NV_NVDLA_CSC_dl_for_check.scala 534:24:@616.4]
  wire [15:0] _T_1219; // @[NV_NVDLA_CSC_dl_for_check.scala 533:24:@617.4]
  wire [15:0] _T_1220; // @[NV_NVDLA_CSC_dl_for_check.scala 532:24:@618.4]
  wire [9:0] _T_1226; // @[NV_NVDLA_CSC_dl_for_check.scala 539:68:@620.4]
  wire [14:0] _T_1227; // @[Cat.scala 30:58:@621.4]
  wire  _T_1238; // @[NV_NVDLA_CSC_dl_for_check.scala 542:68:@632.4]
  wire  _T_1239; // @[NV_NVDLA_CSC_dl_for_check.scala 542:57:@633.4]
  wire  _T_1240; // @[NV_NVDLA_CSC_dl_for_check.scala 542:72:@634.4]
  wire  _T_1241; // @[NV_NVDLA_CSC_dl_for_check.scala 542:88:@635.4]
  wire  _T_1242; // @[NV_NVDLA_CSC_dl_for_check.scala 542:103:@636.4]
  wire  _T_1243; // @[NV_NVDLA_CSC_dl_for_check.scala 542:39:@637.4]
  wire  _T_1245; // @[NV_NVDLA_CSC_dl_for_check.scala 544:42:@639.4]
  wire  _T_1248; // @[NV_NVDLA_CSC_dl_for_check.scala 544:74:@640.4]
  wire  _T_1249; // @[NV_NVDLA_CSC_dl_for_check.scala 544:28:@641.4]
  wire  _T_1251; // @[NV_NVDLA_CSC_dl_for_check.scala 545:36:@643.4]
  wire  _T_1252; // @[NV_NVDLA_CSC_dl_for_check.scala 545:72:@644.4]
  wire  _T_1253; // @[NV_NVDLA_CSC_dl_for_check.scala 545:51:@645.4]
  wire [13:0] _GEN_71; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@646.4]
  wire [15:0] _GEN_72; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@646.4]
  wire [13:0] _GEN_73; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@650.4]
  wire [15:0] _GEN_74; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@650.4]
  wire [15:0] _GEN_75; // @[NV_NVDLA_CSC_dl_for_check.scala 555:26:@654.4]
  reg [13:0] _T_1256; // @[NV_NVDLA_CSC_dl_for_check.scala 561:27:@657.4]
  reg [31:0] _RAND_85;
  reg [13:0] _T_1259; // @[NV_NVDLA_CSC_dl_for_check.scala 562:27:@658.4]
  reg [31:0] _RAND_86;
  wire [13:0] _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@659.4]
  wire [14:0] _T_1261; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@659.4]
  wire [14:0] _T_1262; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@660.4]
  wire [13:0] _T_1263; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@661.4]
  wire [13:0] _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@662.4]
  wire [14:0] _T_1264; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@662.4]
  wire [13:0] _T_1265; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@663.4]
  wire  _T_1266; // @[NV_NVDLA_CSC_dl_for_check.scala 566:52:@664.4]
  wire  _T_1267; // @[NV_NVDLA_CSC_dl_for_check.scala 566:35:@665.4]
  wire [13:0] _T_1270; // @[NV_NVDLA_CSC_dl_for_check.scala 568:25:@668.4]
  wire [13:0] _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 567:25:@669.4]
  wire [13:0] _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 566:25:@670.4]
  wire  _T_1275; // @[NV_NVDLA_CSC_dl_for_check.scala 569:91:@673.4]
  wire  _T_1276; // @[NV_NVDLA_CSC_dl_for_check.scala 569:54:@674.4]
  wire  _T_1277; // @[NV_NVDLA_CSC_dl_for_check.scala 569:36:@675.4]
  wire [5:0] _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@679.4]
  wire [10:0] _T_1281; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@679.4]
  wire [13:0] _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 572:33:@680.4]
  wire [14:0] _T_1282; // @[NV_NVDLA_CSC_dl_for_check.scala 572:33:@680.4]
  wire [13:0] _T_1283; // @[NV_NVDLA_CSC_dl_for_check.scala 572:33:@681.4]
  wire [13:0] _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 572:51:@682.4]
  wire [14:0] _T_1284; // @[NV_NVDLA_CSC_dl_for_check.scala 572:51:@682.4]
  wire [13:0] _T_1285; // @[NV_NVDLA_CSC_dl_for_check.scala 572:51:@683.4]
  wire [13:0] _GEN_76; // @[NV_NVDLA_CSC_dl_for_check.scala 574:26:@684.4]
  wire [13:0] _GEN_77; // @[NV_NVDLA_CSC_dl_for_check.scala 575:26:@687.4]
  wire  _T_1286; // @[NV_NVDLA_CSC_dl_for_check.scala 578:39:@690.4]
  wire [13:0] _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@691.4]
  wire  _T_1287; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@691.4]
  wire  _T_1288; // @[NV_NVDLA_CSC_dl_for_check.scala 578:44:@692.4]
  wire  _T_1289; // @[NV_NVDLA_CSC_dl_for_check.scala 578:92:@693.4]
  wire  _T_1290; // @[NV_NVDLA_CSC_dl_for_check.scala 578:78:@694.4]
  wire [13:0] _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@695.4]
  wire  _T_1291; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@695.4]
  wire  _T_1292; // @[NV_NVDLA_CSC_dl_for_check.scala 578:97:@696.4]
  wire  _T_1305; // @[NV_NVDLA_CSC_dl_for_check.scala 581:42:@706.4]
  wire  _T_1415; // @[NV_NVDLA_CSC_dl_for_check.scala 666:33:@792.4]
  wire  _T_1416; // @[NV_NVDLA_CSC_dl_for_check.scala 667:24:@793.4]
  wire [12:0] _T_1418; // @[NV_NVDLA_CSC_dl_for_check.scala 667:77:@794.4]
  wire [14:0] _T_1419; // @[Cat.scala 30:58:@795.4]
  wire  _T_1421; // @[NV_NVDLA_CSC_dl_for_check.scala 668:38:@796.4]
  wire [11:0] _T_1426; // @[NV_NVDLA_CSC_dl_for_check.scala 669:54:@799.4]
  wire [14:0] _T_1427; // @[Cat.scala 30:58:@800.4]
  wire [14:0] _T_1428; // @[NV_NVDLA_CSC_dl_for_check.scala 668:23:@801.4]
  wire [14:0] _T_1429; // @[NV_NVDLA_CSC_dl_for_check.scala 667:23:@802.4]
  wire [14:0] _T_1430; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@803.4]
  wire [13:0] _T_1431; // @[NV_NVDLA_CSC_dl_for_check.scala 678:24:@805.4]
  wire [11:0] _T_1308; // @[NV_NVDLA_CSC_dl_for_check.scala 585:32:@708.4]
  wire [14:0] _GEN_700; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@709.4]
  wire  _T_1309; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@709.4]
  wire  _T_1310; // @[NV_NVDLA_CSC_dl_for_check.scala 586:34:@710.4]
  wire  _T_1311; // @[NV_NVDLA_CSC_dl_for_check.scala 586:24:@711.4]
  wire  _T_1312; // @[NV_NVDLA_CSC_dl_for_check.scala 587:29:@712.4]
  wire  _T_1313; // @[NV_NVDLA_CSC_dl_for_check.scala 587:33:@713.4]
  wire  _T_1314; // @[NV_NVDLA_CSC_dl_for_check.scala 588:39:@714.4]
  wire  _T_1315; // @[NV_NVDLA_CSC_dl_for_check.scala 588:37:@715.4]
  wire  _T_1316; // @[NV_NVDLA_CSC_dl_for_check.scala 588:56:@716.4]
  wire  _T_1317; // @[NV_NVDLA_CSC_dl_for_check.scala 588:54:@717.4]
  wire  _T_1318; // @[NV_NVDLA_CSC_dl_for_check.scala 591:37:@718.4]
  wire  _T_1319; // @[NV_NVDLA_CSC_dl_for_check.scala 591:27:@719.4]
  wire  _T_1320; // @[NV_NVDLA_CSC_dl_for_check.scala 591:54:@720.4]
  wire  _T_1321; // @[NV_NVDLA_CSC_dl_for_check.scala 591:26:@721.4]
  wire [1:0] _T_1322; // @[NV_NVDLA_CSC_dl_for_check.scala 592:35:@722.4]
  wire  _T_1324; // @[NV_NVDLA_CSC_dl_for_check.scala 593:55:@723.4]
  wire  _T_1325; // @[NV_NVDLA_CSC_dl_for_check.scala 593:42:@724.4]
  wire  _T_1326; // @[NV_NVDLA_CSC_dl_for_check.scala 596:42:@726.4]
  wire [8:0] _T_1330; // @[Cat.scala 30:58:@730.4]
  reg  _T_1333; // @[NV_NVDLA_CSC_dl_for_check.scala 603:31:@731.4]
  reg [31:0] _RAND_87;
  reg [1:0] _T_1336; // @[NV_NVDLA_CSC_dl_for_check.scala 604:31:@732.4]
  reg [31:0] _RAND_88;
  reg [1:0] _T_1339; // @[NV_NVDLA_CSC_dl_for_check.scala 605:31:@733.4]
  reg [31:0] _RAND_89;
  reg  _T_1342; // @[NV_NVDLA_CSC_dl_for_check.scala 606:31:@734.4]
  reg [31:0] _RAND_90;
  reg  _T_1345; // @[NV_NVDLA_CSC_dl_for_check.scala 607:32:@735.4]
  reg [31:0] _RAND_91;
  reg  _T_1348; // @[NV_NVDLA_CSC_dl_for_check.scala 608:31:@736.4]
  reg [31:0] _RAND_92;
  reg [1:0] _T_1351; // @[NV_NVDLA_CSC_dl_for_check.scala 609:35:@737.4]
  reg [31:0] _RAND_93;
  reg  _T_1354; // @[NV_NVDLA_CSC_dl_for_check.scala 610:34:@738.4]
  reg [31:0] _RAND_94;
  reg [8:0] _T_1357; // @[NV_NVDLA_CSC_dl_for_check.scala 611:30:@739.4]
  reg [31:0] _RAND_95;
  reg  _T_1360; // @[NV_NVDLA_CSC_dl_for_check.scala 612:29:@740.4]
  reg [31:0] _RAND_96;
  wire  _T_1361; // @[NV_NVDLA_CSC_dl_for_check.scala 623:38:@750.6]
  wire  _T_1362; // @[NV_NVDLA_CSC_dl_for_check.scala 623:56:@751.6]
  wire [1:0] _GEN_78; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire [1:0] _GEN_79; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_80; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_81; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_82; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire [1:0] _GEN_83; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire [8:0] _GEN_84; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_85; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_86; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_87; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  wire  _GEN_88; // @[NV_NVDLA_CSC_dl_for_check.scala 627:26:@756.4]
  reg [12:0] _T_1365; // @[NV_NVDLA_CSC_dl_for_check.scala 635:21:@759.4]
  reg [31:0] _RAND_97;
  reg [12:0] _T_1368; // @[NV_NVDLA_CSC_dl_for_check.scala 636:24:@760.4]
  reg [31:0] _RAND_98;
  reg [12:0] _T_1371; // @[NV_NVDLA_CSC_dl_for_check.scala 637:26:@761.4]
  reg [31:0] _RAND_99;
  reg [12:0] _T_1374; // @[NV_NVDLA_CSC_dl_for_check.scala 638:26:@762.4]
  reg [31:0] _RAND_100;
  reg [12:0] _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 639:26:@763.4]
  reg [31:0] _RAND_101;
  reg [12:0] _T_1380; // @[NV_NVDLA_CSC_dl_for_check.scala 640:26:@764.4]
  reg [31:0] _RAND_102;
  reg [12:0] _T_1383; // @[NV_NVDLA_CSC_dl_for_check.scala 641:24:@765.4]
  reg [31:0] _RAND_103;
  wire  _T_1384; // @[NV_NVDLA_CSC_dl_for_check.scala 644:32:@766.4]
  wire  _T_1385; // @[NV_NVDLA_CSC_dl_for_check.scala 644:22:@767.4]
  wire [11:0] _T_1386; // @[NV_NVDLA_CSC_dl_for_check.scala 644:49:@768.4]
  wire [11:0] _T_1388; // @[NV_NVDLA_CSC_dl_for_check.scala 644:21:@769.4]
  wire  _T_1390; // @[NV_NVDLA_CSC_dl_for_check.scala 646:34:@770.4]
  wire [12:0] _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@771.4]
  wire [13:0] _T_1392; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@771.4]
  wire [12:0] _T_1393; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@772.4]
  wire [12:0] _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 646:19:@773.4]
  wire [12:0] _T_1395; // @[NV_NVDLA_CSC_dl_for_check.scala 645:19:@774.4]
  wire  _T_1399; // @[NV_NVDLA_CSC_dl_for_check.scala 648:31:@778.4]
  wire [13:0] _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@779.4]
  wire [25:0] _T_1400; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@779.4]
  wire [12:0] _T_1401; // @[NV_NVDLA_CSC_dl_for_check.scala 651:50:@780.4]
  wire [11:0] _GEN_703; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@781.4]
  wire [16:0] _T_1402; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@781.4]
  wire [12:0] _T_1403; // @[NV_NVDLA_CSC_dl_for_check.scala 652:49:@782.4]
  wire [14:0] _GEN_704; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@783.4]
  wire [19:0] _T_1404; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@783.4]
  wire [12:0] _T_1405; // @[NV_NVDLA_CSC_dl_for_check.scala 653:47:@784.4]
  wire [14:0] _GEN_705; // @[NV_NVDLA_CSC_dl_for_check.scala 654:47:@785.4]
  wire [16:0] _T_1407; // @[NV_NVDLA_CSC_dl_for_check.scala 654:47:@785.4]
  wire [16:0] _T_1408; // @[NV_NVDLA_CSC_dl_for_check.scala 654:21:@786.4]
  wire [12:0] _T_1409; // @[NV_NVDLA_CSC_dl_for_check.scala 654:65:@787.4]
  wire  _T_1410; // @[NV_NVDLA_CSC_dl_for_check.scala 655:45:@788.4]
  wire  _T_1411; // @[NV_NVDLA_CSC_dl_for_check.scala 655:34:@789.4]
  wire [1:0] _T_1412; // @[Cat.scala 30:58:@790.4]
  wire [12:0] _GEN_89; // @[NV_NVDLA_CSC_dl_for_check.scala 682:20:@807.4]
  wire [12:0] _GEN_90; // @[NV_NVDLA_CSC_dl_for_check.scala 685:23:@810.4]
  wire  _T_1432; // @[NV_NVDLA_CSC_dl_for_check.scala 688:19:@813.4]
  wire [12:0] _GEN_91; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@814.4]
  wire [12:0] _GEN_92; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@814.4]
  wire [12:0] _GEN_93; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@814.4]
  wire  _T_1433; // @[NV_NVDLA_CSC_dl_for_check.scala 693:19:@819.4]
  wire [12:0] _GEN_94; // @[NV_NVDLA_CSC_dl_for_check.scala 693:23:@820.4]
  wire [13:0] _GEN_95; // @[NV_NVDLA_CSC_dl_for_check.scala 696:20:@823.4]
  reg [12:0] _T_1476_0; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@835.4]
  reg [31:0] _RAND_104;
  reg [12:0] _T_1476_1; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@835.4]
  reg [31:0] _RAND_105;
  reg [12:0] _T_1476_2; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@835.4]
  reg [31:0] _RAND_106;
  reg [12:0] _T_1476_3; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@835.4]
  reg [31:0] _RAND_107;
  reg  _T_1495; // @[NV_NVDLA_CSC_dl_for_check.scala 705:35:@836.4]
  reg [31:0] _RAND_108;
  reg [14:0] _T_1502; // @[NV_NVDLA_CSC_dl_for_check.scala 706:37:@838.4]
  reg [31:0] _RAND_109;
  reg  _T_1505; // @[NV_NVDLA_CSC_dl_for_check.scala 707:32:@839.4]
  reg [31:0] _RAND_110;
  reg [1:0] _T_1511; // @[NV_NVDLA_CSC_dl_for_check.scala 709:33:@841.4]
  reg [31:0] _RAND_111;
  reg [1:0] _T_1514; // @[NV_NVDLA_CSC_dl_for_check.scala 710:33:@842.4]
  reg [31:0] _RAND_112;
  reg  _T_1517; // @[NV_NVDLA_CSC_dl_for_check.scala 711:33:@843.4]
  reg [31:0] _RAND_113;
  reg  _T_1520; // @[NV_NVDLA_CSC_dl_for_check.scala 712:34:@844.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_1523; // @[NV_NVDLA_CSC_dl_for_check.scala 713:33:@845.4]
  reg [31:0] _RAND_115;
  reg  _T_1526; // @[NV_NVDLA_CSC_dl_for_check.scala 714:33:@846.4]
  reg [31:0] _RAND_116;
  reg [1:0] _T_1529; // @[NV_NVDLA_CSC_dl_for_check.scala 715:37:@847.4]
  reg [31:0] _RAND_117;
  reg  _T_1532; // @[NV_NVDLA_CSC_dl_for_check.scala 716:36:@848.4]
  reg [31:0] _RAND_118;
  reg  _T_1535; // @[NV_NVDLA_CSC_dl_for_check.scala 717:31:@849.4]
  reg [31:0] _RAND_119;
  reg [8:0] _T_1538; // @[NV_NVDLA_CSC_dl_for_check.scala 718:32:@850.4]
  reg [31:0] _RAND_120;
  wire [13:0] _T_1539; // @[NV_NVDLA_CSC_dl_for_check.scala 720:29:@851.4]
  wire [12:0] _T_1540; // @[NV_NVDLA_CSC_dl_for_check.scala 720:29:@852.4]
  wire [13:0] _T_1541; // @[NV_NVDLA_CSC_dl_for_check.scala 720:43:@853.4]
  wire [12:0] _T_1542; // @[NV_NVDLA_CSC_dl_for_check.scala 720:43:@854.4]
  wire [13:0] _T_1543; // @[NV_NVDLA_CSC_dl_for_check.scala 720:57:@855.4]
  wire [12:0] _T_1544; // @[NV_NVDLA_CSC_dl_for_check.scala 720:57:@856.4]
  wire [14:0] _GEN_706; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@857.4]
  wire [15:0] _T_1545; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@857.4]
  wire [14:0] _T_1546; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@858.4]
  wire [14:0] _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 721:52:@859.4]
  wire [15:0] _T_1547; // @[NV_NVDLA_CSC_dl_for_check.scala 721:52:@859.4]
  wire [14:0] _T_1548; // @[NV_NVDLA_CSC_dl_for_check.scala 721:52:@860.4]
  wire [14:0] _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 721:64:@861.4]
  wire [15:0] _T_1549; // @[NV_NVDLA_CSC_dl_for_check.scala 721:64:@861.4]
  wire [14:0] _T_1550; // @[NV_NVDLA_CSC_dl_for_check.scala 721:64:@862.4]
  wire  _T_1557; // @[NV_NVDLA_CSC_dl_for_check.scala 722:45:@865.4]
  wire [15:0] _T_1564; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@868.4]
  wire [15:0] _T_1565; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@869.4]
  wire [14:0] _T_1566; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@870.4]
  wire  _T_1567; // @[NV_NVDLA_CSC_dl_for_check.scala 724:35:@871.4]
  wire [14:0] _T_1573; // @[NV_NVDLA_CSC_dl_for_check.scala 725:25:@873.4]
  wire [14:0] _T_1574; // @[NV_NVDLA_CSC_dl_for_check.scala 724:25:@874.4]
  wire  _T_1598; // @[Mux.scala 46:19:@884.4]
  wire [12:0] _T_1599; // @[Mux.scala 46:16:@885.4]
  wire  _T_1600; // @[Mux.scala 46:19:@886.4]
  wire [12:0] _T_1601; // @[Mux.scala 46:16:@887.4]
  wire  _T_1602; // @[Mux.scala 46:19:@888.4]
  wire [12:0] _T_1603; // @[Mux.scala 46:16:@889.4]
  wire  _T_1604; // @[Mux.scala 46:19:@890.4]
  wire [12:0] _T_1605; // @[Mux.scala 46:16:@891.4]
  wire [14:0] _GEN_712; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@892.4]
  wire  _T_1606; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@892.4]
  wire  _T_1607; // @[NV_NVDLA_CSC_dl_for_check.scala 732:85:@893.4]
  wire  _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 732:43:@894.4]
  wire  _T_1609; // @[NV_NVDLA_CSC_dl_for_check.scala 734:38:@895.4]
  wire  _T_1611; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@896.4]
  wire  _T_1612; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@897.4]
  wire  _T_1613; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@898.4]
  wire  _T_1616; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@900.4]
  wire  _T_1617; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@901.4]
  wire  _T_1618; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@902.4]
  wire  _T_1621; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@904.4]
  wire  _T_1622; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@905.4]
  wire  _T_1623; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@906.4]
  wire  _T_1626; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@908.4]
  wire  _T_1627; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@909.4]
  wire  _T_1628; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@910.4]
  wire [14:0] _GEN_96; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@916.4]
  wire [14:0] _GEN_97; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@919.4]
  wire [14:0] _GEN_98; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@922.4]
  wire [14:0] _GEN_99; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@925.4]
  wire  _T_1639; // @[NV_NVDLA_CSC_dl_for_check.scala 747:14:@929.4]
  wire [14:0] _GEN_100; // @[NV_NVDLA_CSC_dl_for_check.scala 747:34:@930.4]
  wire [1:0] _GEN_101; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire [1:0] _GEN_102; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire  _GEN_103; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire  _GEN_104; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire  _GEN_106; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire [1:0] _GEN_107; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire  _GEN_108; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire  _GEN_109; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire [8:0] _GEN_110; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  wire [6:0] _T_1649; // @[Cat.scala 30:58:@957.4]
  wire [28:0] _T_1655; // @[Cat.scala 30:58:@963.4]
  reg  _T_1660; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@965.4]
  reg [31:0] _RAND_121;
  reg  _T_1663; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@966.4]
  reg [31:0] _RAND_122;
  reg  _T_1666; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@967.4]
  reg [31:0] _RAND_123;
  reg  _T_1669; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@968.4]
  reg [31:0] _RAND_124;
  reg  _T_1672; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@969.4]
  reg [31:0] _RAND_125;
  reg  _T_1675; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@970.4]
  reg [31:0] _RAND_126;
  reg [28:0] _T_1680; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@972.4]
  reg [31:0] _RAND_127;
  reg [28:0] _T_1683; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@973.4]
  reg [31:0] _RAND_128;
  reg [28:0] _T_1686; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@974.4]
  reg [31:0] _RAND_129;
  reg [28:0] _T_1689; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@975.4]
  reg [31:0] _RAND_130;
  reg [28:0] _T_1692; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@976.4]
  reg [31:0] _RAND_131;
  reg [28:0] _T_1695; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@977.4]
  reg [31:0] _RAND_132;
  wire [28:0] _GEN_111; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1005.4]
  wire [28:0] _GEN_114; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1014.4]
  wire [28:0] _GEN_117; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1023.4]
  wire [28:0] _GEN_120; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1032.4]
  wire [28:0] _GEN_123; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1041.4]
  wire [28:0] _GEN_126; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1050.4]
  wire [1:0] _T_1756; // @[NV_NVDLA_CSC_dl_for_check.scala 816:41:@1058.4]
  wire [1:0] _T_1757; // @[NV_NVDLA_CSC_dl_for_check.scala 817:41:@1059.4]
  wire  _T_1758; // @[NV_NVDLA_CSC_dl_for_check.scala 818:41:@1060.4]
  wire  _T_1759; // @[NV_NVDLA_CSC_dl_for_check.scala 819:42:@1061.4]
  wire [7:0] _T_1760; // @[NV_NVDLA_CSC_dl_for_check.scala 820:41:@1062.4]
  wire [1:0] _T_1761; // @[NV_NVDLA_CSC_dl_for_check.scala 821:45:@1063.4]
  wire  _T_1764; // @[NV_NVDLA_CSC_dl_for_check.scala 824:39:@1066.4]
  wire [8:0] _T_1765; // @[NV_NVDLA_CSC_dl_for_check.scala 825:40:@1067.4]
  reg  _T_1768; // @[NV_NVDLA_CSC_dl_for_check.scala 830:29:@1068.4]
  reg [31:0] _RAND_133;
  reg  _T_1780; // @[NV_NVDLA_CSC_dl_for_check.scala 834:29:@1072.4]
  reg [31:0] _RAND_134;
  reg [511:0] _T_1791; // @[NV_NVDLA_CSC_dl_for_check.scala 839:19:@1076.4]
  reg [511:0] _RAND_135;
  reg [511:0] _T_1799; // @[NV_NVDLA_CSC_dl_for_check.scala 843:19:@1080.4]
  reg [511:0] _RAND_136;
  wire  _T_1822; // @[NV_NVDLA_CSC_dl_for_check.scala 855:69:@1095.4]
  wire  _T_1823; // @[NV_NVDLA_CSC_dl_for_check.scala 855:74:@1096.4]
  wire  _T_1824; // @[NV_NVDLA_CSC_dl_for_check.scala 855:90:@1097.4]
  wire  _T_1825; // @[NV_NVDLA_CSC_dl_for_check.scala 855:88:@1098.4]
  wire  _T_1865; // @[NV_NVDLA_CSC_dl_for_check.scala 870:22:@1132.4]
  wire  _T_1879; // @[NV_NVDLA_CSC_dl_for_check.scala 874:48:@1143.4]
  wire  _T_1880; // @[NV_NVDLA_CSC_dl_for_check.scala 874:22:@1144.4]
  reg [7:0] _T_1899; // @[NV_NVDLA_CSC_dl_for_check.scala 891:29:@1185.4]
  reg [31:0] _RAND_137;
  reg [7:0] _T_1902; // @[NV_NVDLA_CSC_dl_for_check.scala 892:29:@1186.4]
  reg [31:0] _RAND_138;
  reg [7:0] _T_1905; // @[NV_NVDLA_CSC_dl_for_check.scala 893:29:@1187.4]
  reg [31:0] _RAND_139;
  reg [7:0] _T_1908; // @[NV_NVDLA_CSC_dl_for_check.scala 894:29:@1188.4]
  reg [31:0] _RAND_140;
  reg [7:0] _T_1911; // @[NV_NVDLA_CSC_dl_for_check.scala 895:33:@1189.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_1914; // @[NV_NVDLA_CSC_dl_for_check.scala 896:33:@1190.4]
  reg [31:0] _RAND_142;
  reg [7:0] _T_1917; // @[NV_NVDLA_CSC_dl_for_check.scala 897:33:@1191.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_1920; // @[NV_NVDLA_CSC_dl_for_check.scala 898:33:@1192.4]
  reg [31:0] _RAND_144;
  reg  _T_1931; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1196.4]
  reg [31:0] _RAND_145;
  reg [26:0] _T_1945; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1201.4]
  reg [31:0] _RAND_146;
  wire [26:0] _T_1957; // @[Cat.scala 30:58:@1211.4]
  wire [26:0] _GEN_137; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1214.4]
  wire [26:0] _GEN_138; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1218.4]
  wire [26:0] _GEN_139; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1222.4]
  wire [26:0] _GEN_140; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1226.4]
  wire  _T_1986; // @[NV_NVDLA_CSC_dl_for_check.scala 931:39:@1252.4]
  wire  _T_1987; // @[NV_NVDLA_CSC_dl_for_check.scala 932:39:@1253.4]
  wire  _T_1988; // @[NV_NVDLA_CSC_dl_for_check.scala 933:39:@1254.4]
  wire  _T_1989; // @[NV_NVDLA_CSC_dl_for_check.scala 934:39:@1255.4]
  wire [8:0] _T_1990; // @[NV_NVDLA_CSC_dl_for_check.scala 936:38:@1256.4]
  wire [8:0] _T_1991; // @[NV_NVDLA_CSC_dl_for_check.scala 937:38:@1257.4]
  wire [8:0] _T_1992; // @[NV_NVDLA_CSC_dl_for_check.scala 938:38:@1258.4]
  wire [8:0] _T_1993; // @[NV_NVDLA_CSC_dl_for_check.scala 939:38:@1259.4]
  wire  _T_1994; // @[NV_NVDLA_CSC_dl_for_check.scala 941:44:@1260.4]
  wire  _T_1995; // @[NV_NVDLA_CSC_dl_for_check.scala 942:44:@1261.4]
  wire  _T_1996; // @[NV_NVDLA_CSC_dl_for_check.scala 943:44:@1262.4]
  wire  _T_1997; // @[NV_NVDLA_CSC_dl_for_check.scala 944:44:@1263.4]
  wire [1:0] _T_1998; // @[NV_NVDLA_CSC_dl_for_check.scala 947:31:@1264.4]
  wire [7:0] _T_2002; // @[NV_NVDLA_CSC_dl_for_check.scala 951:31:@1268.4]
  wire [1:0] _T_2003; // @[NV_NVDLA_CSC_dl_for_check.scala 952:35:@1269.4]
  wire [7:0] _T_2013; // @[NV_NVDLA_CSC_dl_for_check.scala 963:29:@1278.4]
  wire  _T_2024; // @[NV_NVDLA_CSC_dl_for_check.scala 968:50:@1282.4]
  wire [7:0] _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1283.4]
  wire [8:0] _T_2026; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1283.4]
  wire [7:0] _T_2027; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1284.4]
  wire [8:0] _T_2028; // @[NV_NVDLA_CSC_dl_for_check.scala 968:133:@1285.4]
  wire [8:0] _T_2029; // @[NV_NVDLA_CSC_dl_for_check.scala 968:133:@1286.4]
  wire [7:0] _T_2030; // @[NV_NVDLA_CSC_dl_for_check.scala 968:133:@1287.4]
  wire [7:0] _T_2031; // @[NV_NVDLA_CSC_dl_for_check.scala 968:29:@1288.4]
  wire [8:0] _T_2035; // @[NV_NVDLA_CSC_dl_for_check.scala 969:111:@1290.4]
  wire [7:0] _T_2036; // @[NV_NVDLA_CSC_dl_for_check.scala 969:111:@1291.4]
  wire [8:0] _T_2037; // @[NV_NVDLA_CSC_dl_for_check.scala 969:133:@1292.4]
  wire [8:0] _T_2038; // @[NV_NVDLA_CSC_dl_for_check.scala 969:133:@1293.4]
  wire [7:0] _T_2039; // @[NV_NVDLA_CSC_dl_for_check.scala 969:133:@1294.4]
  wire [7:0] _T_2040; // @[NV_NVDLA_CSC_dl_for_check.scala 969:29:@1295.4]
  wire [8:0] _T_2044; // @[NV_NVDLA_CSC_dl_for_check.scala 970:111:@1297.4]
  wire [7:0] _T_2045; // @[NV_NVDLA_CSC_dl_for_check.scala 970:111:@1298.4]
  wire [8:0] _T_2046; // @[NV_NVDLA_CSC_dl_for_check.scala 970:133:@1299.4]
  wire [8:0] _T_2047; // @[NV_NVDLA_CSC_dl_for_check.scala 970:133:@1300.4]
  wire [7:0] _T_2048; // @[NV_NVDLA_CSC_dl_for_check.scala 970:133:@1301.4]
  wire [7:0] _T_2049; // @[NV_NVDLA_CSC_dl_for_check.scala 970:29:@1302.4]
  wire [8:0] _T_2053; // @[NV_NVDLA_CSC_dl_for_check.scala 971:111:@1304.4]
  wire [7:0] _T_2054; // @[NV_NVDLA_CSC_dl_for_check.scala 971:111:@1305.4]
  wire [8:0] _T_2055; // @[NV_NVDLA_CSC_dl_for_check.scala 971:133:@1306.4]
  wire [8:0] _T_2056; // @[NV_NVDLA_CSC_dl_for_check.scala 971:133:@1307.4]
  wire [7:0] _T_2057; // @[NV_NVDLA_CSC_dl_for_check.scala 971:133:@1308.4]
  wire [7:0] _T_2058; // @[NV_NVDLA_CSC_dl_for_check.scala 971:29:@1309.4]
  wire  _T_2060; // @[NV_NVDLA_CSC_dl_for_check.scala 980:52:@1310.4]
  wire  _T_2061; // @[NV_NVDLA_CSC_dl_for_check.scala 980:50:@1311.4]
  wire  _T_2062; // @[NV_NVDLA_CSC_dl_for_check.scala 981:50:@1312.4]
  wire [7:0] _T_2067; // @[NV_NVDLA_CSC_dl_for_check.scala 981:27:@1315.4]
  wire [7:0] _T_2068; // @[NV_NVDLA_CSC_dl_for_check.scala 980:27:@1316.4]
  wire [7:0] _T_2069; // @[NV_NVDLA_CSC_dl_for_check.scala 979:27:@1317.4]
  wire  _T_2071; // @[NV_NVDLA_CSC_dl_for_check.scala 985:52:@1318.4]
  wire  _T_2072; // @[NV_NVDLA_CSC_dl_for_check.scala 985:50:@1319.4]
  wire  _T_2073; // @[NV_NVDLA_CSC_dl_for_check.scala 986:50:@1320.4]
  wire [7:0] _T_2078; // @[NV_NVDLA_CSC_dl_for_check.scala 986:27:@1323.4]
  wire [7:0] _T_2079; // @[NV_NVDLA_CSC_dl_for_check.scala 985:27:@1324.4]
  wire [7:0] _T_2080; // @[NV_NVDLA_CSC_dl_for_check.scala 984:27:@1325.4]
  wire  _T_2082; // @[NV_NVDLA_CSC_dl_for_check.scala 990:52:@1326.4]
  wire  _T_2083; // @[NV_NVDLA_CSC_dl_for_check.scala 990:50:@1327.4]
  wire  _T_2084; // @[NV_NVDLA_CSC_dl_for_check.scala 991:50:@1328.4]
  wire [7:0] _T_2089; // @[NV_NVDLA_CSC_dl_for_check.scala 991:27:@1331.4]
  wire [7:0] _T_2090; // @[NV_NVDLA_CSC_dl_for_check.scala 990:27:@1332.4]
  wire [7:0] _T_2091; // @[NV_NVDLA_CSC_dl_for_check.scala 989:27:@1333.4]
  wire  _T_2093; // @[NV_NVDLA_CSC_dl_for_check.scala 995:52:@1334.4]
  wire  _T_2094; // @[NV_NVDLA_CSC_dl_for_check.scala 995:50:@1335.4]
  wire  _T_2095; // @[NV_NVDLA_CSC_dl_for_check.scala 996:50:@1336.4]
  wire [7:0] _T_2100; // @[NV_NVDLA_CSC_dl_for_check.scala 996:27:@1339.4]
  wire [7:0] _T_2101; // @[NV_NVDLA_CSC_dl_for_check.scala 995:27:@1340.4]
  wire [7:0] _T_2102; // @[NV_NVDLA_CSC_dl_for_check.scala 994:27:@1341.4]
  wire  _T_2103; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:46:@1342.4]
  wire  _T_2104; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:51:@1343.4]
  wire  _T_2105; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:34:@1344.4]
  wire  _T_2106; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:46:@1345.4]
  wire  _T_2107; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:51:@1346.4]
  wire  _T_2109; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:87:@1347.4]
  wire  _T_2110; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:69:@1348.4]
  wire  _T_2111; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:34:@1349.4]
  wire  _T_2112; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:46:@1350.4]
  wire  _T_2113; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:51:@1351.4]
  wire  _T_2115; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:87:@1352.4]
  wire  _T_2116; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:69:@1353.4]
  wire  _T_2117; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:34:@1354.4]
  wire  _T_2118; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:46:@1355.4]
  wire  _T_2119; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:51:@1356.4]
  wire  _T_2122; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:69:@1358.4]
  wire  _T_2123; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:34:@1359.4]
  wire  _T_2124; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:50:@1360.4]
  wire  _T_2125; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:55:@1361.4]
  wire  _T_2126; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:73:@1362.4]
  wire  _T_2127; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:97:@1363.4]
  wire  _T_2128; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:38:@1364.4]
  wire  _T_2129; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:50:@1365.4]
  wire  _T_2130; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:55:@1366.4]
  wire  _T_2131; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:73:@1367.4]
  wire  _T_2132; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:97:@1368.4]
  wire  _T_2134; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:138:@1369.4]
  wire  _T_2135; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:120:@1370.4]
  wire  _T_2136; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:38:@1371.4]
  wire  _T_2137; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:50:@1372.4]
  wire  _T_2138; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:55:@1373.4]
  wire  _T_2139; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:73:@1374.4]
  wire  _T_2140; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:97:@1375.4]
  wire  _T_2142; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:138:@1376.4]
  wire  _T_2143; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:120:@1377.4]
  wire  _T_2144; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:38:@1378.4]
  wire  _T_2145; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:50:@1379.4]
  wire  _T_2146; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:55:@1380.4]
  wire  _T_2147; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:73:@1381.4]
  wire  _T_2148; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:97:@1382.4]
  wire  _T_2151; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:120:@1384.4]
  wire  _T_2152; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:38:@1385.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_dl_for_check.scala 1010:24:@1386.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_dl_for_check.scala 1011:24:@1389.4]
  wire [7:0] _GEN_143; // @[NV_NVDLA_CSC_dl_for_check.scala 1012:24:@1392.4]
  wire [7:0] _GEN_144; // @[NV_NVDLA_CSC_dl_for_check.scala 1013:24:@1395.4]
  wire [7:0] _GEN_145; // @[NV_NVDLA_CSC_dl_for_check.scala 1014:28:@1398.4]
  wire [7:0] _GEN_146; // @[NV_NVDLA_CSC_dl_for_check.scala 1015:28:@1401.4]
  wire [7:0] _GEN_147; // @[NV_NVDLA_CSC_dl_for_check.scala 1016:28:@1404.4]
  wire [7:0] _GEN_148; // @[NV_NVDLA_CSC_dl_for_check.scala 1017:28:@1407.4]
  wire [7:0] _T_2153; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:55:@1410.4]
  wire [63:0] _T_2156; // @[Cat.scala 30:58:@1413.4]
  wire [127:0] _T_2157; // @[Cat.scala 30:58:@1414.4]
  wire [255:0] _T_2158; // @[Cat.scala 30:58:@1415.4]
  wire [511:0] _T_2159; // @[Cat.scala 30:58:@1416.4]
  wire [511:0] _T_2160; // @[NV_NVDLA_CSC_dl_for_check.scala 1028:23:@1417.4]
  wire [511:0] _T_2164; // @[NV_NVDLA_CSC_dl_for_check.scala 1033:23:@1421.4]
  wire  _T_2170; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:37:@1426.4]
  wire  _T_2173; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:43:@1427.4]
  wire  _T_2174; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:87:@1428.4]
  wire  _T_2176; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:91:@1429.4]
  wire  _T_2177; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:72:@1430.4]
  wire [255:0] _T_2179; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:171:@1431.4]
  wire [511:0] _T_2180; // @[Cat.scala 30:58:@1432.4]
  wire  _T_2186; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:72:@1436.4]
  wire [255:0] _T_2188; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:171:@1437.4]
  wire [511:0] _T_2189; // @[Cat.scala 30:58:@1438.4]
  wire [511:0] _T_2190; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:27:@1439.4]
  wire [511:0] _T_2191; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:27:@1440.4]
  wire [511:0] _T_2192; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:27:@1441.4]
  wire [7:0] _T_2263; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1444.4]
  wire [7:0] _T_2264; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1446.4]
  wire [7:0] _T_2265; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1448.4]
  wire [7:0] _T_2266; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1450.4]
  wire [7:0] _T_2267; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1452.4]
  wire [7:0] _T_2268; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1454.4]
  wire [7:0] _T_2269; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1456.4]
  wire [7:0] _T_2270; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1458.4]
  wire [7:0] _T_2271; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1460.4]
  wire [7:0] _T_2272; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1462.4]
  wire [7:0] _T_2273; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1464.4]
  wire [7:0] _T_2274; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1466.4]
  wire [7:0] _T_2275; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1468.4]
  wire [7:0] _T_2276; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1470.4]
  wire [7:0] _T_2277; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1472.4]
  wire [7:0] _T_2278; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1474.4]
  wire [7:0] _T_2279; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1476.4]
  wire [7:0] _T_2280; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1478.4]
  wire [7:0] _T_2281; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1480.4]
  wire [7:0] _T_2282; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1482.4]
  wire [7:0] _T_2283; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1484.4]
  wire [7:0] _T_2284; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1486.4]
  wire [7:0] _T_2285; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1488.4]
  wire [7:0] _T_2286; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1490.4]
  wire [7:0] _T_2287; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1492.4]
  wire [7:0] _T_2288; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1494.4]
  wire [7:0] _T_2289; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1496.4]
  wire [7:0] _T_2290; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1498.4]
  wire [7:0] _T_2291; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1500.4]
  wire [7:0] _T_2292; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1502.4]
  wire [7:0] _T_2293; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1504.4]
  wire [7:0] _T_2294; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1506.4]
  wire [7:0] _T_2295; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1508.4]
  wire [7:0] _T_2296; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1510.4]
  wire [7:0] _T_2297; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1512.4]
  wire [7:0] _T_2298; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1514.4]
  wire [7:0] _T_2299; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1516.4]
  wire [7:0] _T_2300; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1518.4]
  wire [7:0] _T_2301; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1520.4]
  wire [7:0] _T_2302; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1522.4]
  wire [7:0] _T_2303; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1524.4]
  wire [7:0] _T_2304; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1526.4]
  wire [7:0] _T_2305; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1528.4]
  wire [7:0] _T_2306; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1530.4]
  wire [7:0] _T_2307; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1532.4]
  wire [7:0] _T_2308; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1534.4]
  wire [7:0] _T_2309; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1536.4]
  wire [7:0] _T_2310; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1538.4]
  wire [7:0] _T_2311; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1540.4]
  wire [7:0] _T_2312; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1542.4]
  wire [7:0] _T_2313; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1544.4]
  wire [7:0] _T_2314; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1546.4]
  wire [7:0] _T_2315; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1548.4]
  wire [7:0] _T_2316; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1550.4]
  wire [7:0] _T_2317; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1552.4]
  wire [7:0] _T_2318; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1554.4]
  wire [7:0] _T_2319; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1556.4]
  wire [7:0] _T_2320; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1558.4]
  wire [7:0] _T_2321; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1560.4]
  wire [7:0] _T_2322; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1562.4]
  wire [7:0] _T_2323; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1564.4]
  wire [7:0] _T_2324; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1566.4]
  wire [7:0] _T_2325; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1568.4]
  wire [7:0] _T_2326; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1570.4]
  reg [255:0] _T_2328; // @[NV_NVDLA_CSC_dl_for_check.scala 1068:28:@1572.4]
  reg [255:0] _RAND_147;
  reg [127:0] _T_2330; // @[NV_NVDLA_CSC_dl_for_check.scala 1069:28:@1573.4]
  reg [127:0] _RAND_148;
  reg [127:0] _T_2332; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:28:@1574.4]
  reg [127:0] _RAND_149;
  reg [127:0] _T_2334; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:28:@1575.4]
  reg [127:0] _RAND_150;
  reg [127:0] _T_2336; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:28:@1576.4]
  reg [127:0] _RAND_151;
  reg [127:0] _T_2338; // @[NV_NVDLA_CSC_dl_for_check.scala 1075:28:@1577.4]
  reg [127:0] _RAND_152;
  wire  _T_2339; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:39:@1578.4]
  wire  _T_2340; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:29:@1579.4]
  wire [1023:0] _T_2342; // @[Cat.scala 30:58:@1580.4]
  wire [1023:0] _T_2343; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:28:@1581.4]
  wire  _T_2344; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:39:@1582.4]
  wire  _T_2345; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:29:@1583.4]
  wire [1023:0] _T_2347; // @[Cat.scala 30:58:@1584.4]
  wire [1023:0] _T_2348; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:28:@1585.4]
  wire  _T_2349; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:39:@1586.4]
  wire  _T_2350; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:29:@1587.4]
  wire [1023:0] _T_2353; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:28:@1589.4]
  wire  _T_2354; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:39:@1590.4]
  wire  _T_2355; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:29:@1591.4]
  wire [1023:0] _T_2358; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:28:@1593.4]
  wire [10:0] _T_2360; // @[Cat.scala 30:58:@1594.4]
  wire [1023:0] _T_2361; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:41:@1595.4]
  wire [511:0] _T_2362; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:82:@1596.4]
  wire [10:0] _T_2364; // @[Cat.scala 30:58:@1597.4]
  wire [1023:0] _T_2365; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:41:@1598.4]
  wire [511:0] _T_2366; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:82:@1599.4]
  wire [10:0] _T_2368; // @[Cat.scala 30:58:@1600.4]
  wire [1023:0] _T_2369; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:41:@1601.4]
  wire [511:0] _T_2370; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:82:@1602.4]
  wire [10:0] _T_2372; // @[Cat.scala 30:58:@1603.4]
  wire [1023:0] _T_2373; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:41:@1604.4]
  wire [511:0] _T_2374; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:82:@1605.4]
  wire  _T_2375; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:36:@1606.4]
  wire  _T_2376; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:26:@1607.4]
  wire  _T_2379; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:41:@1608.4]
  wire [127:0] _T_2380; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:81:@1609.4]
  wire [511:0] _T_2386; // @[Cat.scala 30:58:@1615.4]
  wire  _T_2388; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:41:@1616.4]
  wire [255:0] _T_2389; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:81:@1617.4]
  wire [511:0] _T_2391; // @[Cat.scala 30:58:@1619.4]
  wire [511:0] _T_2393; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:25:@1621.4]
  wire [511:0] _T_2394; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:25:@1622.4]
  wire [511:0] _T_2395; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:25:@1623.4]
  wire [7:0] _T_2466; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1625.4]
  wire [7:0] _T_2467; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1627.4]
  wire [7:0] _T_2468; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1629.4]
  wire [7:0] _T_2469; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1631.4]
  wire [7:0] _T_2470; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1633.4]
  wire [7:0] _T_2471; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1635.4]
  wire [7:0] _T_2472; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1637.4]
  wire [7:0] _T_2473; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1639.4]
  wire [7:0] _T_2474; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1641.4]
  wire [7:0] _T_2475; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1643.4]
  wire [7:0] _T_2476; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1645.4]
  wire [7:0] _T_2477; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1647.4]
  wire [7:0] _T_2478; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1649.4]
  wire [7:0] _T_2479; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1651.4]
  wire [7:0] _T_2480; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1653.4]
  wire [7:0] _T_2481; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1655.4]
  wire [7:0] _T_2482; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1657.4]
  wire [7:0] _T_2483; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1659.4]
  wire [7:0] _T_2484; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1661.4]
  wire [7:0] _T_2485; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1663.4]
  wire [7:0] _T_2486; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1665.4]
  wire [7:0] _T_2487; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1667.4]
  wire [7:0] _T_2488; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1669.4]
  wire [7:0] _T_2489; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1671.4]
  wire [7:0] _T_2490; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1673.4]
  wire [7:0] _T_2491; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1675.4]
  wire [7:0] _T_2492; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1677.4]
  wire [7:0] _T_2493; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1679.4]
  wire [7:0] _T_2494; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1681.4]
  wire [7:0] _T_2495; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1683.4]
  wire [7:0] _T_2496; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1685.4]
  wire [7:0] _T_2497; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1687.4]
  wire [7:0] _T_2498; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1689.4]
  wire [7:0] _T_2499; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1691.4]
  wire [7:0] _T_2500; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1693.4]
  wire [7:0] _T_2501; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1695.4]
  wire [7:0] _T_2502; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1697.4]
  wire [7:0] _T_2503; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1699.4]
  wire [7:0] _T_2504; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1701.4]
  wire [7:0] _T_2505; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1703.4]
  wire [7:0] _T_2506; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1705.4]
  wire [7:0] _T_2507; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1707.4]
  wire [7:0] _T_2508; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1709.4]
  wire [7:0] _T_2509; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1711.4]
  wire [7:0] _T_2510; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1713.4]
  wire [7:0] _T_2511; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1715.4]
  wire [7:0] _T_2512; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1717.4]
  wire [7:0] _T_2513; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1719.4]
  wire [7:0] _T_2514; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1721.4]
  wire [7:0] _T_2515; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1723.4]
  wire [7:0] _T_2516; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1725.4]
  wire [7:0] _T_2517; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1727.4]
  wire [7:0] _T_2518; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1729.4]
  wire [7:0] _T_2519; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1731.4]
  wire [7:0] _T_2520; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1733.4]
  wire [7:0] _T_2521; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1735.4]
  wire [7:0] _T_2522; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1737.4]
  wire [7:0] _T_2523; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1739.4]
  wire [7:0] _T_2524; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1741.4]
  wire [7:0] _T_2525; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1743.4]
  wire [7:0] _T_2526; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1745.4]
  wire [7:0] _T_2527; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1747.4]
  wire [7:0] _T_2528; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1749.4]
  wire [7:0] _T_2529; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1751.4]
  wire  _T_2531; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:59:@1753.4]
  wire  _T_2532; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:41:@1754.4]
  wire  _T_2534; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:59:@1755.4]
  wire  _T_2535; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:41:@1756.4]
  wire  _T_2538; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:41:@1758.4]
  wire [511:0] _GEN_149; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:24:@1759.4]
  wire [255:0] _GEN_150; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1762.4]
  wire [511:0] _GEN_151; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1762.4]
  wire [511:0] _GEN_154; // @[NV_NVDLA_CSC_dl_for_check.scala 1109:24:@1766.4]
  wire [318:0] _T_2544; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:56:@1772.4]
  wire [63:0] _T_2545; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:73:@1773.4]
  wire [63:0] _T_2546; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:24:@1774.4]
  wire  _T_2548; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:51:@1775.4]
  wire [63:0] _T_2555; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:32:@1777.4]
  wire  _T_2557; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:51:@1778.4]
  wire [31:0] _T_2564; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:32:@1780.4]
  wire  _T_2566; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:51:@1781.4]
  wire [31:0] _T_2573; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:32:@1783.4]
  wire [31:0] _T_2574; // @[NV_NVDLA_CSC_dl_for_check.scala 1124:57:@1784.4]
  wire [63:0] _T_2580; // @[Cat.scala 30:58:@1786.4]
  wire [15:0] _T_2581; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:57:@1787.4]
  wire [15:0] _T_2582; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:106:@1788.4]
  wire [15:0] _T_2583; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:155:@1789.4]
  wire [63:0] _T_2591; // @[Cat.scala 30:58:@1793.4]
  wire  _T_2593; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:43:@1794.4]
  wire [15:0] _T_2594; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:89:@1795.4]
  wire [63:0] _T_2596; // @[Cat.scala 30:58:@1797.4]
  wire [63:0] _T_2597; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:116:@1798.4]
  wire  _T_2599; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:43:@1799.4]
  wire [31:0] _T_2600; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:89:@1800.4]
  wire [63:0] _T_2601; // @[Cat.scala 30:58:@1801.4]
  wire [63:0] _T_2602; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:116:@1802.4]
  wire [63:0] _T_2603; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:26:@1803.4]
  wire [63:0] _T_2604; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:26:@1804.4]
  wire  _T_2605; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:35:@1805.4]
  wire [7:0] _T_2606_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire [7:0] _T_2606_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  wire  _T_2739; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1807.4]
  wire  _T_2741; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1808.4]
  wire  _T_2743; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1809.4]
  wire  _T_2745; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1810.4]
  wire  _T_2747; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1811.4]
  wire  _T_2749; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1812.4]
  wire  _T_2751; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1813.4]
  wire  _T_2753; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1814.4]
  wire  _T_2755; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1815.4]
  wire  _T_2757; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1816.4]
  wire  _T_2759; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1817.4]
  wire  _T_2761; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1818.4]
  wire  _T_2763; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1819.4]
  wire  _T_2765; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1820.4]
  wire  _T_2767; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1821.4]
  wire  _T_2769; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1822.4]
  wire  _T_2771; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1823.4]
  wire  _T_2773; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1824.4]
  wire  _T_2775; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1825.4]
  wire  _T_2777; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1826.4]
  wire  _T_2779; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1827.4]
  wire  _T_2781; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1828.4]
  wire  _T_2783; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1829.4]
  wire  _T_2785; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1830.4]
  wire  _T_2787; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1831.4]
  wire  _T_2789; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1832.4]
  wire  _T_2791; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1833.4]
  wire  _T_2793; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1834.4]
  wire  _T_2795; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1835.4]
  wire  _T_2797; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1836.4]
  wire  _T_2799; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1837.4]
  wire  _T_2801; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1838.4]
  wire  _T_2803; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1839.4]
  wire  _T_2805; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1840.4]
  wire  _T_2807; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1841.4]
  wire  _T_2809; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1842.4]
  wire  _T_2811; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1843.4]
  wire  _T_2813; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1844.4]
  wire  _T_2815; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1845.4]
  wire  _T_2817; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1846.4]
  wire  _T_2819; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1847.4]
  wire  _T_2821; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1848.4]
  wire  _T_2823; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1849.4]
  wire  _T_2825; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1850.4]
  wire  _T_2827; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1851.4]
  wire  _T_2829; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1852.4]
  wire  _T_2831; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1853.4]
  wire  _T_2833; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1854.4]
  wire  _T_2835; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1855.4]
  wire  _T_2837; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1856.4]
  wire  _T_2839; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1857.4]
  wire  _T_2841; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1858.4]
  wire  _T_2843; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1859.4]
  wire  _T_2845; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1860.4]
  wire  _T_2847; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1861.4]
  wire  _T_2849; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1862.4]
  wire  _T_2851; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1863.4]
  wire  _T_2853; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1864.4]
  wire  _T_2855; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1865.4]
  wire  _T_2857; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1866.4]
  wire  _T_2859; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1867.4]
  wire  _T_2861; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1868.4]
  wire  _T_2863; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1869.4]
  wire  _T_2865; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1870.4]
  wire  _T_2936; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1936.4]
  wire  _T_2937; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1937.4]
  wire  _T_2938; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1938.4]
  wire  _T_2939; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1939.4]
  wire  _T_2940; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1940.4]
  wire  _T_2941; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1941.4]
  wire  _T_2942; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1942.4]
  wire  _T_2943; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1943.4]
  wire  _T_2944; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1944.4]
  wire  _T_2945; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1945.4]
  wire  _T_2946; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1946.4]
  wire  _T_2947; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1947.4]
  wire  _T_2948; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1948.4]
  wire  _T_2949; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1949.4]
  wire  _T_2950; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1950.4]
  wire  _T_2951; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1951.4]
  wire  _T_2952; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1952.4]
  wire  _T_2953; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1953.4]
  wire  _T_2954; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1954.4]
  wire  _T_2955; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1955.4]
  wire  _T_2956; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1956.4]
  wire  _T_2957; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1957.4]
  wire  _T_2958; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1958.4]
  wire  _T_2959; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1959.4]
  wire  _T_2960; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1960.4]
  wire  _T_2961; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1961.4]
  wire  _T_2962; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1962.4]
  wire  _T_2963; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1963.4]
  wire  _T_2964; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1964.4]
  wire  _T_2965; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1965.4]
  wire  _T_2966; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1966.4]
  wire  _T_2967; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1967.4]
  wire  _T_2968; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1968.4]
  wire  _T_2969; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1969.4]
  wire  _T_2970; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1970.4]
  wire  _T_2971; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1971.4]
  wire  _T_2972; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1972.4]
  wire  _T_2973; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1973.4]
  wire  _T_2974; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1974.4]
  wire  _T_2975; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1975.4]
  wire  _T_2976; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1976.4]
  wire  _T_2977; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1977.4]
  wire  _T_2978; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1978.4]
  wire  _T_2979; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1979.4]
  wire  _T_2980; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1980.4]
  wire  _T_2981; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1981.4]
  wire  _T_2982; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1982.4]
  wire  _T_2983; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1983.4]
  wire  _T_2984; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1984.4]
  wire  _T_2985; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1985.4]
  wire  _T_2986; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1986.4]
  wire  _T_2987; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1987.4]
  wire  _T_2988; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1988.4]
  wire  _T_2989; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1989.4]
  wire  _T_2990; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1990.4]
  wire  _T_2991; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1991.4]
  wire  _T_2992; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1992.4]
  wire  _T_2993; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1993.4]
  wire  _T_2994; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1994.4]
  wire  _T_2995; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1995.4]
  wire  _T_2996; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1996.4]
  wire  _T_2997; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1997.4]
  wire  _T_2998; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1998.4]
  wire  _T_2999; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1999.4]
  wire  _T_3000; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2000.4]
  wire  _T_3001; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2001.4]
  wire  _T_3002; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2002.4]
  wire  _T_3003; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2003.4]
  wire  _T_3004; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2004.4]
  wire  _T_3005; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2005.4]
  wire  _T_3006; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2006.4]
  wire  _T_3007; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2007.4]
  wire  _T_3008; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2008.4]
  wire  _T_3009; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2009.4]
  wire  _T_3010; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2010.4]
  wire  _T_3011; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2011.4]
  wire  _T_3012; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2012.4]
  wire  _T_3013; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2013.4]
  wire  _T_3014; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2014.4]
  wire  _T_3015; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2015.4]
  wire  _T_3016; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2016.4]
  wire  _T_3017; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2017.4]
  wire  _T_3018; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2018.4]
  wire  _T_3019; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2019.4]
  wire  _T_3020; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2020.4]
  wire  _T_3021; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2021.4]
  wire  _T_3022; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2022.4]
  wire  _T_3023; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2023.4]
  wire  _T_3024; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2024.4]
  wire  _T_3025; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2025.4]
  wire  _T_3026; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2026.4]
  wire  _T_3027; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2027.4]
  wire  _T_3028; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2028.4]
  wire  _T_3029; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2029.4]
  wire  _T_3030; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2030.4]
  wire  _T_3031; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2031.4]
  wire  _T_3032; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2032.4]
  wire  _T_3033; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2033.4]
  wire  _T_3034; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2034.4]
  wire  _T_3035; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2035.4]
  wire  _T_3036; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2036.4]
  wire  _T_3037; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2037.4]
  wire  _T_3038; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2038.4]
  wire  _T_3039; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2039.4]
  wire  _T_3040; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2040.4]
  wire  _T_3041; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2041.4]
  wire  _T_3042; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2042.4]
  wire  _T_3043; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2043.4]
  wire  _T_3044; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2044.4]
  wire  _T_3045; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2045.4]
  wire  _T_3046; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2046.4]
  wire  _T_3047; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2047.4]
  wire  _T_3048; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2048.4]
  wire  _T_3049; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2049.4]
  wire  _T_3050; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2050.4]
  wire  _T_3051; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2051.4]
  wire  _T_3052; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2052.4]
  wire  _T_3053; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2053.4]
  wire  _T_3054; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2054.4]
  wire  _T_3055; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2055.4]
  wire  _T_3056; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2056.4]
  wire  _T_3057; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2057.4]
  wire  _T_3058; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2058.4]
  wire  _T_3059; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2059.4]
  wire  _T_3060; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2060.4]
  wire  _T_3061; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2061.4]
  wire  _T_3062; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2062.4]
  wire  _T_3063; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2063.4]
  reg  _T_3136; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:27:@2129.4]
  reg [31:0] _RAND_153;
  reg  _T_3406_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_154;
  reg  _T_3406_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_155;
  reg  _T_3406_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_156;
  reg  _T_3406_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_157;
  reg  _T_3406_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_158;
  reg  _T_3406_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_159;
  reg  _T_3406_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_160;
  reg  _T_3406_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_161;
  reg  _T_3406_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_162;
  reg  _T_3406_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_163;
  reg  _T_3406_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_164;
  reg  _T_3406_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_165;
  reg  _T_3406_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_166;
  reg  _T_3406_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_167;
  reg  _T_3406_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_168;
  reg  _T_3406_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_169;
  reg  _T_3406_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_170;
  reg  _T_3406_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_171;
  reg  _T_3406_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_172;
  reg  _T_3406_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_173;
  reg  _T_3406_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_174;
  reg  _T_3406_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_175;
  reg  _T_3406_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_176;
  reg  _T_3406_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_177;
  reg  _T_3406_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_178;
  reg  _T_3406_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_179;
  reg  _T_3406_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_180;
  reg  _T_3406_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_181;
  reg  _T_3406_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_182;
  reg  _T_3406_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_183;
  reg  _T_3406_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_184;
  reg  _T_3406_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_185;
  reg  _T_3406_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_186;
  reg  _T_3406_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_187;
  reg  _T_3406_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_188;
  reg  _T_3406_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_189;
  reg  _T_3406_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_190;
  reg  _T_3406_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_191;
  reg  _T_3406_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_192;
  reg  _T_3406_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_193;
  reg  _T_3406_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_194;
  reg  _T_3406_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_195;
  reg  _T_3406_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_196;
  reg  _T_3406_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_197;
  reg  _T_3406_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_198;
  reg  _T_3406_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_199;
  reg  _T_3406_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_200;
  reg  _T_3406_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_201;
  reg  _T_3406_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_202;
  reg  _T_3406_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_203;
  reg  _T_3406_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_204;
  reg  _T_3406_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_205;
  reg  _T_3406_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_206;
  reg  _T_3406_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_207;
  reg  _T_3406_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_208;
  reg  _T_3406_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_209;
  reg  _T_3406_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_210;
  reg  _T_3406_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_211;
  reg  _T_3406_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_212;
  reg  _T_3406_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_213;
  reg  _T_3406_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_214;
  reg  _T_3406_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_215;
  reg  _T_3406_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_216;
  reg  _T_3406_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2196.4]
  reg [31:0] _RAND_217;
  reg [7:0] _T_3606_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_218;
  reg [7:0] _T_3606_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_219;
  reg [7:0] _T_3606_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_220;
  reg [7:0] _T_3606_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_221;
  reg [7:0] _T_3606_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_222;
  reg [7:0] _T_3606_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_223;
  reg [7:0] _T_3606_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_224;
  reg [7:0] _T_3606_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_225;
  reg [7:0] _T_3606_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_226;
  reg [7:0] _T_3606_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_227;
  reg [7:0] _T_3606_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_228;
  reg [7:0] _T_3606_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_229;
  reg [7:0] _T_3606_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_230;
  reg [7:0] _T_3606_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_231;
  reg [7:0] _T_3606_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_232;
  reg [7:0] _T_3606_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_233;
  reg [7:0] _T_3606_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_234;
  reg [7:0] _T_3606_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_235;
  reg [7:0] _T_3606_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_236;
  reg [7:0] _T_3606_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_237;
  reg [7:0] _T_3606_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_238;
  reg [7:0] _T_3606_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_239;
  reg [7:0] _T_3606_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_240;
  reg [7:0] _T_3606_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_241;
  reg [7:0] _T_3606_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_242;
  reg [7:0] _T_3606_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_243;
  reg [7:0] _T_3606_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_244;
  reg [7:0] _T_3606_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_245;
  reg [7:0] _T_3606_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_246;
  reg [7:0] _T_3606_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_247;
  reg [7:0] _T_3606_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_248;
  reg [7:0] _T_3606_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_249;
  reg [7:0] _T_3606_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_250;
  reg [7:0] _T_3606_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_251;
  reg [7:0] _T_3606_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_252;
  reg [7:0] _T_3606_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_253;
  reg [7:0] _T_3606_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_254;
  reg [7:0] _T_3606_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_255;
  reg [7:0] _T_3606_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_256;
  reg [7:0] _T_3606_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_3606_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_3606_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_3606_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_3606_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_3606_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_3606_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_3606_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_3606_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_3606_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_3606_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_3606_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_3606_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_3606_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_3606_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_3606_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_3606_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_3606_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_3606_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_3606_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_3606_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_3606_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_3606_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_3606_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_3606_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2197.4]
  reg [31:0] _RAND_281;
  wire  _GEN_156; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_209; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  wire  _T_3673; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2268.4]
  wire  _T_3674; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2272.4]
  wire  _T_3675; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2276.4]
  wire  _T_3676; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2280.4]
  wire  _T_3677; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2284.4]
  wire  _T_3678; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2288.4]
  wire  _T_3679; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2292.4]
  wire  _T_3680; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2296.4]
  wire  _T_3681; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2300.4]
  wire  _T_3682; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2304.4]
  wire  _T_3683; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2308.4]
  wire  _T_3684; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2312.4]
  wire  _T_3685; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2316.4]
  wire  _T_3686; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2320.4]
  wire  _T_3687; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2324.4]
  wire  _T_3688; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2328.4]
  wire  _T_3689; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2332.4]
  wire  _T_3690; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2336.4]
  wire  _T_3691; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2340.4]
  wire  _T_3692; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2344.4]
  wire  _T_3693; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2348.4]
  wire  _T_3694; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2352.4]
  wire  _T_3695; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2356.4]
  wire  _T_3696; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2360.4]
  wire  _T_3697; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2364.4]
  wire  _T_3698; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2368.4]
  wire  _T_3699; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2372.4]
  wire  _T_3700; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2376.4]
  wire  _T_3701; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2380.4]
  wire  _T_3702; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2384.4]
  wire  _T_3703; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2388.4]
  wire  _T_3704; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2392.4]
  wire  _T_3705; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2396.4]
  wire  _T_3706; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2400.4]
  wire  _T_3707; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2404.4]
  wire  _T_3708; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2408.4]
  wire  _T_3709; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2412.4]
  wire  _T_3710; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2416.4]
  wire  _T_3711; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2420.4]
  wire  _T_3712; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2424.4]
  wire  _T_3713; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2428.4]
  wire  _T_3714; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2432.4]
  wire  _T_3715; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2436.4]
  wire  _T_3716; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2440.4]
  wire  _T_3717; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2444.4]
  wire  _T_3718; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2448.4]
  wire  _T_3719; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2452.4]
  wire  _T_3720; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2456.4]
  wire  _T_3721; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2460.4]
  wire  _T_3722; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2464.4]
  wire  _T_3723; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2468.4]
  wire  _T_3724; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2472.4]
  wire  _T_3725; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2476.4]
  wire  _T_3726; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2480.4]
  wire  _T_3727; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2484.4]
  wire  _T_3728; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2488.4]
  wire  _T_3729; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2492.4]
  wire  _T_3730; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2496.4]
  wire  _T_3731; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2500.4]
  wire  _T_3732; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2504.4]
  wire  _T_3733; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2508.4]
  wire  _T_3734; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2512.4]
  wire  _T_3735; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2516.4]
  wire  _T_3736; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2520.4]
  reg  _T_3739; // @[NV_NVDLA_CSC_dl_for_check.scala 1169:26:@2524.4]
  reg [31:0] _RAND_282;
  reg  _T_4006_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_283;
  reg  _T_4006_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_284;
  reg  _T_4006_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_285;
  reg  _T_4006_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_286;
  reg  _T_4006_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_287;
  reg  _T_4006_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_288;
  reg  _T_4006_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_289;
  reg  _T_4006_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_290;
  reg  _T_4006_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_291;
  reg  _T_4006_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_292;
  reg  _T_4006_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_293;
  reg  _T_4006_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_294;
  reg  _T_4006_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_295;
  reg  _T_4006_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_296;
  reg  _T_4006_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_297;
  reg  _T_4006_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_298;
  reg  _T_4006_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_299;
  reg  _T_4006_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_300;
  reg  _T_4006_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_301;
  reg  _T_4006_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_302;
  reg  _T_4006_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_303;
  reg  _T_4006_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_304;
  reg  _T_4006_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_305;
  reg  _T_4006_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_306;
  reg  _T_4006_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_307;
  reg  _T_4006_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_308;
  reg  _T_4006_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_309;
  reg  _T_4006_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_310;
  reg  _T_4006_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_311;
  reg  _T_4006_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_312;
  reg  _T_4006_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_313;
  reg  _T_4006_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_314;
  reg  _T_4006_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_315;
  reg  _T_4006_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_316;
  reg  _T_4006_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_317;
  reg  _T_4006_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_318;
  reg  _T_4006_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_319;
  reg  _T_4006_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_320;
  reg  _T_4006_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_321;
  reg  _T_4006_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_322;
  reg  _T_4006_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_323;
  reg  _T_4006_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_324;
  reg  _T_4006_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_325;
  reg  _T_4006_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_326;
  reg  _T_4006_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_327;
  reg  _T_4006_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_328;
  reg  _T_4006_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_329;
  reg  _T_4006_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_330;
  reg  _T_4006_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_331;
  reg  _T_4006_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_332;
  reg  _T_4006_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_333;
  reg  _T_4006_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_334;
  reg  _T_4006_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_335;
  reg  _T_4006_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_336;
  reg  _T_4006_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_337;
  reg  _T_4006_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_338;
  reg  _T_4006_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_339;
  reg  _T_4006_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_340;
  reg  _T_4006_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_341;
  reg  _T_4006_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_342;
  reg  _T_4006_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_343;
  reg  _T_4006_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_344;
  reg  _T_4006_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_345;
  reg  _T_4006_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2590.4]
  reg [31:0] _RAND_346;
  reg [8:0] _T_4205; // @[NV_NVDLA_CSC_dl_for_check.scala 1171:26:@2591.4]
  reg [31:0] _RAND_347;
  reg [7:0] _T_4209_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_348;
  reg [7:0] _T_4209_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_349;
  reg [7:0] _T_4209_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_350;
  reg [7:0] _T_4209_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_351;
  reg [7:0] _T_4209_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_352;
  reg [7:0] _T_4209_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_353;
  reg [7:0] _T_4209_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_354;
  reg [7:0] _T_4209_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_355;
  reg [7:0] _T_4209_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_356;
  reg [7:0] _T_4209_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_357;
  reg [7:0] _T_4209_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_358;
  reg [7:0] _T_4209_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_359;
  reg [7:0] _T_4209_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_360;
  reg [7:0] _T_4209_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_361;
  reg [7:0] _T_4209_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_362;
  reg [7:0] _T_4209_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_363;
  reg [7:0] _T_4209_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_364;
  reg [7:0] _T_4209_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_365;
  reg [7:0] _T_4209_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_366;
  reg [7:0] _T_4209_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_367;
  reg [7:0] _T_4209_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_368;
  reg [7:0] _T_4209_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_369;
  reg [7:0] _T_4209_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_370;
  reg [7:0] _T_4209_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_371;
  reg [7:0] _T_4209_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_372;
  reg [7:0] _T_4209_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_373;
  reg [7:0] _T_4209_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_374;
  reg [7:0] _T_4209_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_375;
  reg [7:0] _T_4209_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_376;
  reg [7:0] _T_4209_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_377;
  reg [7:0] _T_4209_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_378;
  reg [7:0] _T_4209_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_379;
  reg [7:0] _T_4209_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_380;
  reg [7:0] _T_4209_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_381;
  reg [7:0] _T_4209_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_382;
  reg [7:0] _T_4209_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_383;
  reg [7:0] _T_4209_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_384;
  reg [7:0] _T_4209_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_385;
  reg [7:0] _T_4209_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_386;
  reg [7:0] _T_4209_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_387;
  reg [7:0] _T_4209_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_388;
  reg [7:0] _T_4209_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_389;
  reg [7:0] _T_4209_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_390;
  reg [7:0] _T_4209_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_391;
  reg [7:0] _T_4209_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_392;
  reg [7:0] _T_4209_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_393;
  reg [7:0] _T_4209_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_394;
  reg [7:0] _T_4209_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_395;
  reg [7:0] _T_4209_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_396;
  reg [7:0] _T_4209_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_397;
  reg [7:0] _T_4209_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_398;
  reg [7:0] _T_4209_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_399;
  reg [7:0] _T_4209_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_400;
  reg [7:0] _T_4209_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_401;
  reg [7:0] _T_4209_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_402;
  reg [7:0] _T_4209_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_403;
  reg [7:0] _T_4209_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_404;
  reg [7:0] _T_4209_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_405;
  reg [7:0] _T_4209_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_406;
  reg [7:0] _T_4209_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_407;
  reg [7:0] _T_4209_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_408;
  reg [7:0] _T_4209_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_409;
  reg [7:0] _T_4209_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_410;
  reg [7:0] _T_4209_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2592.4]
  reg [31:0] _RAND_411;
  wire  _T_4276; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:24:@2593.4]
  wire  _T_4411_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4411_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  wire  _T_4543; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:19:@2661.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_289; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  wire [8:0] _GEN_348; // @[NV_NVDLA_CSC_dl_for_check.scala 1182:19:@2728.4]
  reg  _T_4546; // @[NV_NVDLA_CSC_dl_for_check.scala 1195:29:@2923.4]
  reg [31:0] _RAND_412;
  wire  _T_4547; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:27:@2925.4]
  wire [8:0] _T_4549; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:26:@2926.4]
  reg  _T_4552; // @[NV_NVDLA_CSC_dl_for_check.scala 1198:33:@2927.4]
  reg [31:0] _RAND_413;
  reg  _T_4555; // @[NV_NVDLA_CSC_dl_for_check.scala 1199:33:@2930.4]
  reg [31:0] _RAND_414;
  wire  _T_4557; // @[NV_NVDLA_CSC_dl_for_check.scala 1200:85:@2933.4]
  reg [8:0] _T_4559; // @[Reg.scala 19:20:@2934.4]
  reg [31:0] _RAND_415;
  wire [8:0] _GEN_413; // @[Reg.scala 20:19:@2935.4]
  reg [8:0] _T_4563; // @[Reg.scala 19:20:@2940.4]
  reg [31:0] _RAND_416;
  wire [8:0] _GEN_414; // @[Reg.scala 20:19:@2941.4]
  reg  _T_4831_0; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_417;
  reg  _T_4831_1; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_418;
  reg  _T_4831_2; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_419;
  reg  _T_4831_3; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_420;
  reg  _T_4831_4; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_421;
  reg  _T_4831_5; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_422;
  reg  _T_4831_6; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_423;
  reg  _T_4831_7; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_424;
  reg  _T_4831_8; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_425;
  reg  _T_4831_9; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_426;
  reg  _T_4831_10; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_427;
  reg  _T_4831_11; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_428;
  reg  _T_4831_12; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_429;
  reg  _T_4831_13; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_430;
  reg  _T_4831_14; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_431;
  reg  _T_4831_15; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_432;
  reg  _T_4831_16; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_433;
  reg  _T_4831_17; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_434;
  reg  _T_4831_18; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_435;
  reg  _T_4831_19; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_436;
  reg  _T_4831_20; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_437;
  reg  _T_4831_21; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_438;
  reg  _T_4831_22; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_439;
  reg  _T_4831_23; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_440;
  reg  _T_4831_24; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_441;
  reg  _T_4831_25; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_442;
  reg  _T_4831_26; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_443;
  reg  _T_4831_27; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_444;
  reg  _T_4831_28; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_445;
  reg  _T_4831_29; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_446;
  reg  _T_4831_30; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_447;
  reg  _T_4831_31; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_448;
  reg  _T_4831_32; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_449;
  reg  _T_4831_33; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_450;
  reg  _T_4831_34; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_451;
  reg  _T_4831_35; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_452;
  reg  _T_4831_36; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_453;
  reg  _T_4831_37; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_454;
  reg  _T_4831_38; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_455;
  reg  _T_4831_39; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_456;
  reg  _T_4831_40; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_457;
  reg  _T_4831_41; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_458;
  reg  _T_4831_42; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_459;
  reg  _T_4831_43; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_460;
  reg  _T_4831_44; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_461;
  reg  _T_4831_45; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_462;
  reg  _T_4831_46; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_463;
  reg  _T_4831_47; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_464;
  reg  _T_4831_48; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_465;
  reg  _T_4831_49; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_466;
  reg  _T_4831_50; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_467;
  reg  _T_4831_51; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_468;
  reg  _T_4831_52; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_469;
  reg  _T_4831_53; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_470;
  reg  _T_4831_54; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_471;
  reg  _T_4831_55; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_472;
  reg  _T_4831_56; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_473;
  reg  _T_4831_57; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_474;
  reg  _T_4831_58; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_475;
  reg  _T_4831_59; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_476;
  reg  _T_4831_60; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_477;
  reg  _T_4831_61; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_478;
  reg  _T_4831_62; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_479;
  reg  _T_4831_63; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_480;
  wire  _GEN_415; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_416; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_417; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_418; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_419; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_420; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_421; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_422; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_423; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_424; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_425; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_426; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_427; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_428; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_429; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_430; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_431; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_432; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_433; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_434; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_435; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_436; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_437; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_438; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_439; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_440; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_441; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_442; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_443; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_444; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_445; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_446; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_447; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_448; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_449; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_450; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_451; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_452; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_453; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_454; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_455; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_456; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_457; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_458; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_459; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_460; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_461; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_462; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_463; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_464; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_465; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_466; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_467; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_468; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_469; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_470; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_471; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_472; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_473; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_474; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_475; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_476; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_477; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_478; // @[Reg.scala 20:19:@3012.4]
  wire [7:0] _T_5034; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3084.4]
  wire [15:0] _T_5042; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3092.4]
  wire [7:0] _T_5049; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3099.4]
  wire [31:0] _T_5058; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3108.4]
  wire [7:0] _T_5065; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3115.4]
  wire [15:0] _T_5073; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3123.4]
  wire [7:0] _T_5080; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3130.4]
  wire [31:0] _T_5089; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3139.4]
  reg  _T_5358_0; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_481;
  reg  _T_5358_1; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_482;
  reg  _T_5358_2; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_483;
  reg  _T_5358_3; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_484;
  reg  _T_5358_4; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_485;
  reg  _T_5358_5; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_486;
  reg  _T_5358_6; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_487;
  reg  _T_5358_7; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_488;
  reg  _T_5358_8; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_489;
  reg  _T_5358_9; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_490;
  reg  _T_5358_10; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_491;
  reg  _T_5358_11; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_492;
  reg  _T_5358_12; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_493;
  reg  _T_5358_13; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_494;
  reg  _T_5358_14; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_495;
  reg  _T_5358_15; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_496;
  reg  _T_5358_16; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_497;
  reg  _T_5358_17; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_498;
  reg  _T_5358_18; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_499;
  reg  _T_5358_19; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_500;
  reg  _T_5358_20; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_501;
  reg  _T_5358_21; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_502;
  reg  _T_5358_22; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_503;
  reg  _T_5358_23; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_504;
  reg  _T_5358_24; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_505;
  reg  _T_5358_25; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_506;
  reg  _T_5358_26; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_507;
  reg  _T_5358_27; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_508;
  reg  _T_5358_28; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_509;
  reg  _T_5358_29; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_510;
  reg  _T_5358_30; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_511;
  reg  _T_5358_31; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_512;
  reg  _T_5358_32; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_513;
  reg  _T_5358_33; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_514;
  reg  _T_5358_34; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_515;
  reg  _T_5358_35; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_516;
  reg  _T_5358_36; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_517;
  reg  _T_5358_37; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_518;
  reg  _T_5358_38; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_519;
  reg  _T_5358_39; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_520;
  reg  _T_5358_40; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_521;
  reg  _T_5358_41; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_522;
  reg  _T_5358_42; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_523;
  reg  _T_5358_43; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_524;
  reg  _T_5358_44; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_525;
  reg  _T_5358_45; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_526;
  reg  _T_5358_46; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_527;
  reg  _T_5358_47; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_528;
  reg  _T_5358_48; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_529;
  reg  _T_5358_49; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_530;
  reg  _T_5358_50; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_531;
  reg  _T_5358_51; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_532;
  reg  _T_5358_52; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_533;
  reg  _T_5358_53; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_534;
  reg  _T_5358_54; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_535;
  reg  _T_5358_55; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_536;
  reg  _T_5358_56; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_537;
  reg  _T_5358_57; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_538;
  reg  _T_5358_58; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_539;
  reg  _T_5358_59; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_540;
  reg  _T_5358_60; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_541;
  reg  _T_5358_61; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_542;
  reg  _T_5358_62; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_543;
  reg  _T_5358_63; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_544;
  wire  _GEN_479; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_480; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_481; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_482; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_483; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_484; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_485; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_486; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_487; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_488; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_489; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_490; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_491; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_492; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_493; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_494; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_495; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_496; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_497; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_498; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_499; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_500; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_501; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_502; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_503; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_504; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_505; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_506; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_507; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_508; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_509; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_510; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_511; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_512; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_513; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_514; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_515; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_516; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_517; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_518; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_519; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_520; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_521; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_522; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_523; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_524; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_525; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_526; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_527; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_528; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_529; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_530; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_531; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_532; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_533; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_534; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_535; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_536; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_537; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_538; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_539; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_540; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_541; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_542; // @[Reg.scala 20:19:@3209.4]
  wire [7:0] _T_5561; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3281.4]
  wire [15:0] _T_5569; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3289.4]
  wire [7:0] _T_5576; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3296.4]
  wire [31:0] _T_5585; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3305.4]
  wire [7:0] _T_5592; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3312.4]
  wire [15:0] _T_5600; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3320.4]
  wire [7:0] _T_5607; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3327.4]
  wire [31:0] _T_5616; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3336.4]
  reg [7:0] _T_5619; // @[Reg.scala 11:16:@3339.4]
  reg [31:0] _RAND_545;
  reg [7:0] _T_5621; // @[Reg.scala 11:16:@3344.4]
  reg [31:0] _RAND_546;
  reg [7:0] _T_5623; // @[Reg.scala 11:16:@3349.4]
  reg [31:0] _RAND_547;
  reg [7:0] _T_5625; // @[Reg.scala 11:16:@3354.4]
  reg [31:0] _RAND_548;
  reg [7:0] _T_5627; // @[Reg.scala 11:16:@3359.4]
  reg [31:0] _RAND_549;
  reg [7:0] _T_5629; // @[Reg.scala 11:16:@3364.4]
  reg [31:0] _RAND_550;
  reg [7:0] _T_5631; // @[Reg.scala 11:16:@3369.4]
  reg [31:0] _RAND_551;
  reg [7:0] _T_5633; // @[Reg.scala 11:16:@3374.4]
  reg [31:0] _RAND_552;
  reg [7:0] _T_5635; // @[Reg.scala 11:16:@3379.4]
  reg [31:0] _RAND_553;
  reg [7:0] _T_5637; // @[Reg.scala 11:16:@3384.4]
  reg [31:0] _RAND_554;
  reg [7:0] _T_5639; // @[Reg.scala 11:16:@3389.4]
  reg [31:0] _RAND_555;
  reg [7:0] _T_5641; // @[Reg.scala 11:16:@3394.4]
  reg [31:0] _RAND_556;
  reg [7:0] _T_5643; // @[Reg.scala 11:16:@3399.4]
  reg [31:0] _RAND_557;
  reg [7:0] _T_5645; // @[Reg.scala 11:16:@3404.4]
  reg [31:0] _RAND_558;
  reg [7:0] _T_5647; // @[Reg.scala 11:16:@3409.4]
  reg [31:0] _RAND_559;
  reg [7:0] _T_5649; // @[Reg.scala 11:16:@3414.4]
  reg [31:0] _RAND_560;
  reg [7:0] _T_5651; // @[Reg.scala 11:16:@3419.4]
  reg [31:0] _RAND_561;
  reg [7:0] _T_5653; // @[Reg.scala 11:16:@3424.4]
  reg [31:0] _RAND_562;
  reg [7:0] _T_5655; // @[Reg.scala 11:16:@3429.4]
  reg [31:0] _RAND_563;
  reg [7:0] _T_5657; // @[Reg.scala 11:16:@3434.4]
  reg [31:0] _RAND_564;
  reg [7:0] _T_5659; // @[Reg.scala 11:16:@3439.4]
  reg [31:0] _RAND_565;
  reg [7:0] _T_5661; // @[Reg.scala 11:16:@3444.4]
  reg [31:0] _RAND_566;
  reg [7:0] _T_5663; // @[Reg.scala 11:16:@3449.4]
  reg [31:0] _RAND_567;
  reg [7:0] _T_5665; // @[Reg.scala 11:16:@3454.4]
  reg [31:0] _RAND_568;
  reg [7:0] _T_5667; // @[Reg.scala 11:16:@3459.4]
  reg [31:0] _RAND_569;
  reg [7:0] _T_5669; // @[Reg.scala 11:16:@3464.4]
  reg [31:0] _RAND_570;
  reg [7:0] _T_5671; // @[Reg.scala 11:16:@3469.4]
  reg [31:0] _RAND_571;
  reg [7:0] _T_5673; // @[Reg.scala 11:16:@3474.4]
  reg [31:0] _RAND_572;
  reg [7:0] _T_5675; // @[Reg.scala 11:16:@3479.4]
  reg [31:0] _RAND_573;
  reg [7:0] _T_5677; // @[Reg.scala 11:16:@3484.4]
  reg [31:0] _RAND_574;
  reg [7:0] _T_5679; // @[Reg.scala 11:16:@3489.4]
  reg [31:0] _RAND_575;
  reg [7:0] _T_5681; // @[Reg.scala 11:16:@3494.4]
  reg [31:0] _RAND_576;
  reg [7:0] _T_5683; // @[Reg.scala 11:16:@3499.4]
  reg [31:0] _RAND_577;
  reg [7:0] _T_5685; // @[Reg.scala 11:16:@3504.4]
  reg [31:0] _RAND_578;
  reg [7:0] _T_5687; // @[Reg.scala 11:16:@3509.4]
  reg [31:0] _RAND_579;
  reg [7:0] _T_5689; // @[Reg.scala 11:16:@3514.4]
  reg [31:0] _RAND_580;
  reg [7:0] _T_5691; // @[Reg.scala 11:16:@3519.4]
  reg [31:0] _RAND_581;
  reg [7:0] _T_5693; // @[Reg.scala 11:16:@3524.4]
  reg [31:0] _RAND_582;
  reg [7:0] _T_5695; // @[Reg.scala 11:16:@3529.4]
  reg [31:0] _RAND_583;
  reg [7:0] _T_5697; // @[Reg.scala 11:16:@3534.4]
  reg [31:0] _RAND_584;
  reg [7:0] _T_5699; // @[Reg.scala 11:16:@3539.4]
  reg [31:0] _RAND_585;
  reg [7:0] _T_5701; // @[Reg.scala 11:16:@3544.4]
  reg [31:0] _RAND_586;
  reg [7:0] _T_5703; // @[Reg.scala 11:16:@3549.4]
  reg [31:0] _RAND_587;
  reg [7:0] _T_5705; // @[Reg.scala 11:16:@3554.4]
  reg [31:0] _RAND_588;
  reg [7:0] _T_5707; // @[Reg.scala 11:16:@3559.4]
  reg [31:0] _RAND_589;
  reg [7:0] _T_5709; // @[Reg.scala 11:16:@3564.4]
  reg [31:0] _RAND_590;
  reg [7:0] _T_5711; // @[Reg.scala 11:16:@3569.4]
  reg [31:0] _RAND_591;
  reg [7:0] _T_5713; // @[Reg.scala 11:16:@3574.4]
  reg [31:0] _RAND_592;
  reg [7:0] _T_5715; // @[Reg.scala 11:16:@3579.4]
  reg [31:0] _RAND_593;
  reg [7:0] _T_5717; // @[Reg.scala 11:16:@3584.4]
  reg [31:0] _RAND_594;
  reg [7:0] _T_5719; // @[Reg.scala 11:16:@3589.4]
  reg [31:0] _RAND_595;
  reg [7:0] _T_5721; // @[Reg.scala 11:16:@3594.4]
  reg [31:0] _RAND_596;
  reg [7:0] _T_5723; // @[Reg.scala 11:16:@3599.4]
  reg [31:0] _RAND_597;
  reg [7:0] _T_5725; // @[Reg.scala 11:16:@3604.4]
  reg [31:0] _RAND_598;
  reg [7:0] _T_5727; // @[Reg.scala 11:16:@3609.4]
  reg [31:0] _RAND_599;
  reg [7:0] _T_5729; // @[Reg.scala 11:16:@3614.4]
  reg [31:0] _RAND_600;
  reg [7:0] _T_5731; // @[Reg.scala 11:16:@3619.4]
  reg [31:0] _RAND_601;
  reg [7:0] _T_5733; // @[Reg.scala 11:16:@3624.4]
  reg [31:0] _RAND_602;
  reg [7:0] _T_5735; // @[Reg.scala 11:16:@3629.4]
  reg [31:0] _RAND_603;
  reg [7:0] _T_5737; // @[Reg.scala 11:16:@3634.4]
  reg [31:0] _RAND_604;
  reg [7:0] _T_5739; // @[Reg.scala 11:16:@3639.4]
  reg [31:0] _RAND_605;
  reg [7:0] _T_5741; // @[Reg.scala 11:16:@3644.4]
  reg [31:0] _RAND_606;
  reg [7:0] _T_5743; // @[Reg.scala 11:16:@3649.4]
  reg [31:0] _RAND_607;
  reg [7:0] _T_5745; // @[Reg.scala 11:16:@3654.4]
  reg [31:0] _RAND_608;
  reg [7:0] _T_5747; // @[Reg.scala 11:16:@3659.4]
  reg [31:0] _RAND_609;
  reg [7:0] _T_5749; // @[Reg.scala 11:16:@3664.4]
  reg [31:0] _RAND_610;
  reg [7:0] _T_5751; // @[Reg.scala 11:16:@3669.4]
  reg [31:0] _RAND_611;
  reg [7:0] _T_5753; // @[Reg.scala 11:16:@3674.4]
  reg [31:0] _RAND_612;
  reg [7:0] _T_5755; // @[Reg.scala 11:16:@3679.4]
  reg [31:0] _RAND_613;
  reg [7:0] _T_5757; // @[Reg.scala 11:16:@3684.4]
  reg [31:0] _RAND_614;
  reg [7:0] _T_5759; // @[Reg.scala 11:16:@3689.4]
  reg [31:0] _RAND_615;
  reg [7:0] _T_5761; // @[Reg.scala 11:16:@3694.4]
  reg [31:0] _RAND_616;
  reg [7:0] _T_5763; // @[Reg.scala 11:16:@3699.4]
  reg [31:0] _RAND_617;
  reg [7:0] _T_5765; // @[Reg.scala 11:16:@3704.4]
  reg [31:0] _RAND_618;
  reg [7:0] _T_5767; // @[Reg.scala 11:16:@3709.4]
  reg [31:0] _RAND_619;
  reg [7:0] _T_5769; // @[Reg.scala 11:16:@3714.4]
  reg [31:0] _RAND_620;
  reg [7:0] _T_5771; // @[Reg.scala 11:16:@3719.4]
  reg [31:0] _RAND_621;
  reg [7:0] _T_5773; // @[Reg.scala 11:16:@3724.4]
  reg [31:0] _RAND_622;
  reg [7:0] _T_5775; // @[Reg.scala 11:16:@3729.4]
  reg [31:0] _RAND_623;
  reg [7:0] _T_5777; // @[Reg.scala 11:16:@3734.4]
  reg [31:0] _RAND_624;
  reg [7:0] _T_5779; // @[Reg.scala 11:16:@3739.4]
  reg [31:0] _RAND_625;
  reg [7:0] _T_5781; // @[Reg.scala 11:16:@3744.4]
  reg [31:0] _RAND_626;
  reg [7:0] _T_5783; // @[Reg.scala 11:16:@3749.4]
  reg [31:0] _RAND_627;
  reg [7:0] _T_5785; // @[Reg.scala 11:16:@3754.4]
  reg [31:0] _RAND_628;
  reg [7:0] _T_5787; // @[Reg.scala 11:16:@3759.4]
  reg [31:0] _RAND_629;
  reg [7:0] _T_5789; // @[Reg.scala 11:16:@3764.4]
  reg [31:0] _RAND_630;
  reg [7:0] _T_5791; // @[Reg.scala 11:16:@3769.4]
  reg [31:0] _RAND_631;
  reg [7:0] _T_5793; // @[Reg.scala 11:16:@3774.4]
  reg [31:0] _RAND_632;
  reg [7:0] _T_5795; // @[Reg.scala 11:16:@3779.4]
  reg [31:0] _RAND_633;
  reg [7:0] _T_5797; // @[Reg.scala 11:16:@3784.4]
  reg [31:0] _RAND_634;
  reg [7:0] _T_5799; // @[Reg.scala 11:16:@3789.4]
  reg [31:0] _RAND_635;
  reg [7:0] _T_5801; // @[Reg.scala 11:16:@3794.4]
  reg [31:0] _RAND_636;
  reg [7:0] _T_5803; // @[Reg.scala 11:16:@3799.4]
  reg [31:0] _RAND_637;
  reg [7:0] _T_5805; // @[Reg.scala 11:16:@3804.4]
  reg [31:0] _RAND_638;
  reg [7:0] _T_5807; // @[Reg.scala 11:16:@3809.4]
  reg [31:0] _RAND_639;
  reg [7:0] _T_5809; // @[Reg.scala 11:16:@3814.4]
  reg [31:0] _RAND_640;
  reg [7:0] _T_5811; // @[Reg.scala 11:16:@3819.4]
  reg [31:0] _RAND_641;
  reg [7:0] _T_5813; // @[Reg.scala 11:16:@3824.4]
  reg [31:0] _RAND_642;
  reg [7:0] _T_5815; // @[Reg.scala 11:16:@3829.4]
  reg [31:0] _RAND_643;
  reg [7:0] _T_5817; // @[Reg.scala 11:16:@3834.4]
  reg [31:0] _RAND_644;
  reg [7:0] _T_5819; // @[Reg.scala 11:16:@3839.4]
  reg [31:0] _RAND_645;
  reg [7:0] _T_5821; // @[Reg.scala 11:16:@3844.4]
  reg [31:0] _RAND_646;
  reg [7:0] _T_5823; // @[Reg.scala 11:16:@3849.4]
  reg [31:0] _RAND_647;
  reg [7:0] _T_5825; // @[Reg.scala 11:16:@3854.4]
  reg [31:0] _RAND_648;
  reg [7:0] _T_5827; // @[Reg.scala 11:16:@3859.4]
  reg [31:0] _RAND_649;
  reg [7:0] _T_5829; // @[Reg.scala 11:16:@3864.4]
  reg [31:0] _RAND_650;
  reg [7:0] _T_5831; // @[Reg.scala 11:16:@3869.4]
  reg [31:0] _RAND_651;
  reg [7:0] _T_5833; // @[Reg.scala 11:16:@3874.4]
  reg [31:0] _RAND_652;
  reg [7:0] _T_5835; // @[Reg.scala 11:16:@3879.4]
  reg [31:0] _RAND_653;
  reg [7:0] _T_5837; // @[Reg.scala 11:16:@3884.4]
  reg [31:0] _RAND_654;
  reg [7:0] _T_5839; // @[Reg.scala 11:16:@3889.4]
  reg [31:0] _RAND_655;
  reg [7:0] _T_5841; // @[Reg.scala 11:16:@3894.4]
  reg [31:0] _RAND_656;
  reg [7:0] _T_5843; // @[Reg.scala 11:16:@3899.4]
  reg [31:0] _RAND_657;
  reg [7:0] _T_5845; // @[Reg.scala 11:16:@3904.4]
  reg [31:0] _RAND_658;
  reg [7:0] _T_5847; // @[Reg.scala 11:16:@3909.4]
  reg [31:0] _RAND_659;
  reg [7:0] _T_5849; // @[Reg.scala 11:16:@3914.4]
  reg [31:0] _RAND_660;
  reg [7:0] _T_5851; // @[Reg.scala 11:16:@3919.4]
  reg [31:0] _RAND_661;
  reg [7:0] _T_5853; // @[Reg.scala 11:16:@3924.4]
  reg [31:0] _RAND_662;
  reg [7:0] _T_5855; // @[Reg.scala 11:16:@3929.4]
  reg [31:0] _RAND_663;
  reg [7:0] _T_5857; // @[Reg.scala 11:16:@3934.4]
  reg [31:0] _RAND_664;
  reg [7:0] _T_5859; // @[Reg.scala 11:16:@3939.4]
  reg [31:0] _RAND_665;
  reg [7:0] _T_5861; // @[Reg.scala 11:16:@3944.4]
  reg [31:0] _RAND_666;
  reg [7:0] _T_5863; // @[Reg.scala 11:16:@3949.4]
  reg [31:0] _RAND_667;
  reg [7:0] _T_5865; // @[Reg.scala 11:16:@3954.4]
  reg [31:0] _RAND_668;
  reg [7:0] _T_5867; // @[Reg.scala 11:16:@3959.4]
  reg [31:0] _RAND_669;
  reg [7:0] _T_5869; // @[Reg.scala 11:16:@3964.4]
  reg [31:0] _RAND_670;
  reg [7:0] _T_5871; // @[Reg.scala 11:16:@3969.4]
  reg [31:0] _RAND_671;
  reg [7:0] _T_5873; // @[Reg.scala 11:16:@3974.4]
  reg [31:0] _RAND_672;
  assign _T_337 = nvdla_core_rstn == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 95:38:@8.4]
  assign _T_339 = sc_state == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 99:31:@9.4]
  assign _T_343 = sc_state == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 101:31:@11.4]
  assign _T_347 = reg2dp_op_en & _T_339; // @[NV_NVDLA_CSC_dl_for_check.scala 108:32:@14.4]
  assign _T_351 = reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 110:35:@16.4]
  assign _T_352 = _T_351 & reg2dp_datain_format; // @[NV_NVDLA_CSC_dl_for_check.scala 111:22:@17.4]
  assign _T_357 = 7'h9 << reg2dp_y_extension; // @[NV_NVDLA_CSC_dl_for_check.scala 118:53:@18.4]
  assign _T_359 = _T_352 ? _T_357 : 7'h8; // @[NV_NVDLA_CSC_dl_for_check.scala 118:24:@19.4]
  assign _T_360 = _T_359[5:3]; // @[NV_NVDLA_CSC_dl_for_check.scala 118:100:@20.4]
  assign _T_362 = _T_352 ? _T_360 : 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 119:22:@21.4]
  assign _T_364 = _T_362 - 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@22.4]
  assign _T_365 = $unsigned(_T_364); // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@23.4]
  assign _T_367 = reg2dp_conv_x_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 121:51:@24.4]
  assign _T_368 = reg2dp_datain_channel_ext[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 122:62:@25.4]
  assign _T_371 = {_T_367,2'h0}; // @[Cat.scala 30:58:@26.4]
  assign _T_374 = {_T_367,1'h0}; // @[Cat.scala 30:58:@27.4]
  assign _GEN_671 = {{1'd0}, _T_367}; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  assign _T_375 = _T_374 + _GEN_671; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  assign _T_376 = 2'h2 == _T_368; // @[Mux.scala 46:19:@29.4]
  assign _T_377 = _T_376 ? _T_375 : {{2'd0}, _T_367}; // @[Mux.scala 46:16:@30.4]
  assign _T_378 = 2'h3 == _T_368; // @[Mux.scala 46:19:@31.4]
  assign _T_379 = _T_378 ? _T_371 : _T_377; // @[Mux.scala 46:16:@32.4]
  assign _T_381 = reg2dp_weight_channel_ext >= 13'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 126:88:@33.4]
  assign _T_387 = reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 126:172:@35.4]
  assign _T_388 = _T_381 ? 6'h3f : _T_387; // @[NV_NVDLA_CSC_dl_for_check.scala 126:58:@36.4]
  assign _T_391 = {_T_379,1'h0}; // @[Cat.scala 30:58:@37.4]
  assign _GEN_672 = {{1'd0}, _T_379}; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  assign _T_392 = _T_391 + _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  assign _T_393 = _T_391 + _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@39.4]
  assign _GEN_673 = {{1'd0}, _T_387}; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  assign _T_395 = _T_393 + _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  assign _T_396 = _T_393 + _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@42.4]
  assign _T_399 = _T_379 + _T_387; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@44.4]
  assign _T_400 = _T_379 + _T_387; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@45.4]
  assign _T_401 = 2'h1 == reg2dp_y_extension; // @[Mux.scala 46:19:@46.4]
  assign _T_402 = _T_401 ? _T_400 : _T_388; // @[Mux.scala 46:16:@47.4]
  assign _T_403 = 2'h2 == reg2dp_y_extension; // @[Mux.scala 46:19:@48.4]
  assign _T_404 = _T_403 ? _T_396 : {{1'd0}, _T_402}; // @[Mux.scala 46:16:@49.4]
  assign _T_407 = _T_387 + 6'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 129:80:@51.4]
  assign _T_410 = {_T_379,2'h0}; // @[Cat.scala 30:58:@52.4]
  assign _T_415 = _T_401 ? _T_391 : {{1'd0}, _T_379}; // @[Mux.scala 46:16:@55.4]
  assign _T_417 = _T_403 ? _T_410 : {{1'd0}, _T_415}; // @[Mux.scala 46:16:@57.4]
  assign _T_419 = {_T_379,6'h0}; // @[Cat.scala 30:58:@58.4]
  assign _T_421 = reg2dp_conv_y_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 139:52:@59.4]
  assign _T_424 = reg2dp_x_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 140:60:@60.4]
  assign _T_425 = _T_352 ? 6'h1 : _T_424; // @[NV_NVDLA_CSC_dl_for_check.scala 140:21:@61.4]
  assign _T_428 = reg2dp_y_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 141:60:@62.4]
  assign _T_429 = _T_352 ? 6'h1 : _T_428; // @[NV_NVDLA_CSC_dl_for_check.scala 141:21:@63.4]
  assign _T_511 = reg2dp_entries + 14'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 157:43:@87.4]
  assign _T_513 = _T_511 * 15'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 158:41:@89.4]
  assign _T_514 = _T_513[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 158:56:@90.4]
  assign _T_515 = 6'h1 * _T_429; // @[NV_NVDLA_CSC_dl_for_check.scala 160:37:@91.4]
  assign _GEN_674 = {{9'd0}, _T_439}; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  assign _T_516 = _T_460 * _GEN_674; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  assign _T_517 = _T_516[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 161:47:@93.4]
  assign _GEN_675 = {{1'd0}, _T_453}; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  assign _T_518 = _T_460 * _GEN_675; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  assign _T_519 = _T_518[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 162:51:@95.4]
  assign _T_521 = reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 163:41:@96.4]
  assign _T_522 = reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 163:41:@97.4]
  assign _T_524 = reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 164:77:@98.4]
  assign _GEN_676 = {{1'd0}, reg2dp_rls_slices}; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@99.4]
  assign _T_525 = reg2dp_datain_height_ext - _GEN_676; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@99.4]
  assign _T_526 = $unsigned(_T_525); // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@100.4]
  assign _T_527 = reg2dp_skip_data_rls ? _T_524 : _T_526; // @[NV_NVDLA_CSC_dl_for_check.scala 164:23:@101.4]
  assign _T_528 = _T_432 ? _T_446 : _T_509; // @[NV_NVDLA_CSC_dl_for_check.scala 165:24:@102.4]
  assign _GEN_677 = {{1'd0}, _T_528}; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@103.4]
  assign _T_529 = _T_467 * _GEN_677; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@103.4]
  assign _T_530 = _T_529[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 166:54:@104.4]
  assign _T_755 = _T_352 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@175.6]
  assign _T_757 = reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@177.6]
  assign _T_758 = reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@178.6]
  assign _T_760 = reg2dp_datain_width_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 216:48:@180.6]
  assign _T_766 = reg2dp_weight_channel_ext[12:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 219:93:@185.6]
  assign _T_767 = {4'h0,_T_766}; // @[Cat.scala 30:58:@186.6]
  assign _T_771 = {1'h0,reg2dp_entries}; // @[Cat.scala 30:58:@219.6]
  assign _GEN_1 = _T_347 ? _T_755 : _T_548; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_2 = _T_347 ? _T_758 : _T_555; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_3 = _T_347 ? _T_760 : _T_562; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_4 = _T_347 ? reg2dp_datain_width_ext : _T_569; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_5 = _T_347 ? reg2dp_datain_height_ext : _T_576; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_6 = _T_347 ? _T_767 : _T_583; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_7 = _T_347 ? _T_360 : _T_586; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_8 = _T_347 ? _T_360 : _T_589; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_10 = _T_347 ? _T_360 : _T_595; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_11 = _T_347 ? _T_360 : _T_598; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_12 = _T_347 ? _T_360 : _T_601; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_13 = _T_347 ? _T_360 : _T_604; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_15 = _T_347 ? _T_360 : _T_610; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_16 = _T_347 ? _T_360 : _T_613; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_18 = _T_347 ? _T_360 : _T_619; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_19 = _T_347 ? _T_362 : _T_622; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_20 = _T_347 ? _T_362 : _T_625; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_21 = _T_347 ? _T_367 : _T_632; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_22 = _T_347 ? _T_421 : _T_639; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_24 = _T_347 ? 6'h1 : _T_439; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_25 = _T_347 ? 5'h0 : _T_649; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_26 = _T_347 ? _T_404 : _T_656; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_27 = _T_347 ? _T_407 : _T_663; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_28 = _T_347 ? _T_417 : _T_670; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_29 = _T_347 ? {{1'd0}, _T_379} : _T_677; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_30 = _T_347 ? _T_419 : _T_684; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_31 = _T_347 ? _T_425 : _T_691; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_32 = _T_347 ? _T_429 : _T_698; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_33 = _T_347 ? reg2dp_pad_value : _T_705; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_34 = _T_347 ? _T_511 : _T_460; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_35 = _T_347 ? _T_514 : _T_467; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_36 = _T_347 ? _T_771 : _T_712; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_37 = _T_347 ? {{2'd0}, _T_515} : _T_453; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_38 = _T_347 ? {{2'd0}, _T_522} : _T_446; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_39 = _T_347 ? _T_527 : _T_509; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_40 = _T_347 ? reg2dp_dataout_width : _T_474; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@171.4]
  assign _GEN_43 = _T_432 ? _T_517 : _T_495; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  assign _GEN_44 = _T_432 ? _T_519 : _T_502; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  assign _GEN_45 = _T_432 ? _T_460 : _T_719; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  assign _GEN_46 = _T_432 ? _T_460 : _T_726; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  assign _GEN_47 = _T_432 ? _T_530 : _T_488; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@232.4]
  assign _GEN_48 = _T_343 ? _T_509 : _T_733; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@239.4]
  assign _GEN_49 = _T_343 ? _T_530 : _T_740; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@239.4]
  assign _T_873 = _T_733 != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 328:37:@314.4]
  assign _T_874 = sg2dl_reuse_rls & _T_873; // @[NV_NVDLA_CSC_dl_for_check.scala 328:23:@315.4]
  assign _T_1958 = _T_595[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 918:32:@1229.4]
  assign _T_1959 = _T_1958 & _T_1934; // @[NV_NVDLA_CSC_dl_for_check.scala 918:36:@1230.4]
  assign _T_1960 = _T_595[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 919:35:@1231.4]
  assign _T_1961 = _T_1960 & _T_1928; // @[NV_NVDLA_CSC_dl_for_check.scala 919:39:@1232.4]
  assign _T_1962 = _T_1959 | _T_1961; // @[NV_NVDLA_CSC_dl_for_check.scala 918:57:@1233.4]
  assign _T_1963 = _T_595[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 920:35:@1234.4]
  assign _T_1964 = _T_1963 & _T_1925; // @[NV_NVDLA_CSC_dl_for_check.scala 920:39:@1235.4]
  assign _T_1965 = _T_1962 | _T_1964; // @[NV_NVDLA_CSC_dl_for_check.scala 919:60:@1236.4]
  assign _T_1966 = _T_598[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 927:42:@1238.4]
  assign _T_1970 = _T_1966 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1240.4]
  assign _T_1971 = _T_1970 & _T_1948; // @[NV_NVDLA_CSC_dl_for_check.scala 927:47:@1241.4]
  assign _T_1972 = _T_598[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 928:42:@1242.4]
  assign _T_1976 = _T_1972 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1244.4]
  assign _T_1977 = _T_1976 & _T_1942; // @[NV_NVDLA_CSC_dl_for_check.scala 928:47:@1245.4]
  assign _T_1978 = _T_1971 | _T_1977; // @[NV_NVDLA_CSC_dl_for_check.scala 927:66:@1246.4]
  assign _T_1979 = _T_598[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 929:42:@1247.4]
  assign _T_1983 = _T_1979 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1249.4]
  assign _T_1984 = _T_1983 & _T_1939; // @[NV_NVDLA_CSC_dl_for_check.scala 929:47:@1250.4]
  assign _T_1985 = _T_1978 | _T_1984; // @[NV_NVDLA_CSC_dl_for_check.scala 928:66:@1251.4]
  assign _T_2004 = _T_1985[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 953:26:@1270.4]
  assign _T_871 = _T_1965 & _T_2004; // @[NV_NVDLA_CSC_dl_for_check.scala 325:29:@313.4]
  assign _T_876 = _T_446 != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 328:66:@316.4]
  assign _T_877 = _T_871 & _T_876; // @[NV_NVDLA_CSC_dl_for_check.scala 328:53:@317.4]
  assign _T_878 = _T_874 | _T_877; // @[NV_NVDLA_CSC_dl_for_check.scala 328:42:@318.4]
  assign _T_879 = _T_871 ? _T_446 : _T_733; // @[NV_NVDLA_CSC_dl_for_check.scala 329:28:@320.4]
  assign _T_880 = _T_871 ? _T_488 : _T_740; // @[NV_NVDLA_CSC_dl_for_check.scala 330:29:@322.4]
  assign _T_811 = _T_878 ? _T_880 : 15'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 297:28:@262.4]
  assign _T_819 = _T_793 + _T_811; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@269.4]
  assign _T_820 = _T_793 + _T_811; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@270.4]
  assign _T_826 = {_T_555,9'h0}; // @[Cat.scala 30:58:@272.4]
  assign _GEN_678 = {{1'd0}, _T_826}; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@273.4]
  assign _T_827 = _T_820 - _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@273.4]
  assign _T_828 = $unsigned(_T_827); // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@274.4]
  assign _T_829 = _T_828[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@275.4]
  assign _T_836 = _T_820 >= _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 304:45:@278.4]
  assign _T_838 = _T_836 ? _T_829 : _T_820; // @[NV_NVDLA_CSC_dl_for_check.scala 305:83:@279.4]
  assign _T_839 = sc2cdma_dat_pending_req ? 15'h0 : _T_838; // @[NV_NVDLA_CSC_dl_for_check.scala 305:25:@280.4]
  assign _T_865 = _T_878 | sc2cdma_dat_pending_req; // @[NV_NVDLA_CSC_dl_for_check.scala 316:13:@303.4]
  assign _GEN_52 = _T_865 ? _T_839 : _T_793; // @[NV_NVDLA_CSC_dl_for_check.scala 316:25:@304.4]
  assign _GEN_54 = _T_878 ? _T_879 : _T_886; // @[Reg.scala 20:19:@328.4]
  assign _GEN_55 = _T_878 ? _T_880 : _T_889; // @[Reg.scala 20:19:@333.4]
  assign _T_939 = {{30'd0}, _T_906}; // @[NV_NVDLA_CSC_dl_for_check.scala 365:19:@376.4 NV_NVDLA_CSC_dl_for_check.scala 369:12:@382.4]
  assign _GEN_61 = _T_906 ? _T_939 : _T_942; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@384.4]
  assign _GEN_62 = _T_928 ? _T_942 : _T_945; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@388.4]
  assign _GEN_63 = _T_931 ? _T_945 : _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@392.4]
  assign _GEN_64 = _T_934 ? _T_948 : _T_951; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@396.4]
  assign _T_952 = _T_586[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 378:30:@399.4]
  assign _T_953 = _T_952 & _T_928; // @[NV_NVDLA_CSC_dl_for_check.scala 378:34:@400.4]
  assign _T_954 = _T_586[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 379:30:@401.4]
  assign _T_955 = _T_954 & _T_934; // @[NV_NVDLA_CSC_dl_for_check.scala 379:34:@402.4]
  assign _T_956 = _T_953 | _T_955; // @[NV_NVDLA_CSC_dl_for_check.scala 378:50:@403.4]
  assign _T_957 = _T_586[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 380:30:@404.4]
  assign _T_958 = _T_957 & _T_937; // @[NV_NVDLA_CSC_dl_for_check.scala 380:34:@405.4]
  assign _T_959 = _T_956 | _T_958; // @[NV_NVDLA_CSC_dl_for_check.scala 379:50:@406.4]
  assign _T_960 = _T_589[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 382:37:@407.4]
  assign _T_964 = _T_960 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@409.4]
  assign _T_965 = _T_964 & _T_942; // @[NV_NVDLA_CSC_dl_for_check.scala 382:42:@410.4]
  assign _T_966 = _T_589[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 383:37:@411.4]
  assign _T_970 = _T_966 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@413.4]
  assign _T_971 = _T_970 & _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 383:42:@414.4]
  assign _T_972 = _T_965 | _T_971; // @[NV_NVDLA_CSC_dl_for_check.scala 382:56:@415.4]
  assign _T_973 = _T_589[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 384:37:@416.4]
  assign _T_977 = _T_973 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@418.4]
  assign _T_978 = _T_977 & _T_951; // @[NV_NVDLA_CSC_dl_for_check.scala 384:42:@419.4]
  assign _T_979 = _T_972 | _T_978; // @[NV_NVDLA_CSC_dl_for_check.scala 383:56:@420.4]
  assign _T_980 = _T_979[4:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 387:24:@421.4]
  assign _T_981 = _T_979[9:5]; // @[NV_NVDLA_CSC_dl_for_check.scala 388:24:@422.4]
  assign _T_982 = _T_979[16:10]; // @[NV_NVDLA_CSC_dl_for_check.scala 389:28:@423.4]
  assign _T_983 = _T_979[23:17]; // @[NV_NVDLA_CSC_dl_for_check.scala 390:29:@424.4]
  assign _T_984 = _T_979[25:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 391:25:@425.4]
  assign _T_985 = _T_979[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 392:25:@426.4]
  assign _T_986 = _T_979[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 393:27:@427.4]
  assign _T_987 = _T_979[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 394:25:@428.4]
  assign _T_988 = _T_979[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 395:25:@429.4]
  assign _T_989 = _T_979[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 396:27:@430.4]
  assign _T_1000 = _T_996 + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 405:24:@434.4]
  assign _T_1001 = _T_996 + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 405:24:@435.4]
  assign _T_1004 = _T_996 == _T_649; // @[NV_NVDLA_CSC_dl_for_check.scala 407:27:@439.4]
  assign _T_1002 = _T_1004 ? 5'h0 : _T_1001; // @[NV_NVDLA_CSC_dl_for_check.scala 404:17:@436.4]
  assign _T_1003 = _T_347 ? 5'h0 : _T_1002; // @[NV_NVDLA_CSC_dl_for_check.scala 403:17:@437.4]
  assign _T_1011 = _T_1007 + 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 413:31:@443.4]
  assign _T_1012 = _T_1007 + 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 413:31:@444.4]
  assign _GEN_682 = {{1'd0}, _T_1012}; // @[NV_NVDLA_CSC_dl_for_check.scala 414:32:@445.4]
  assign _T_1013 = _GEN_682 == _T_622; // @[NV_NVDLA_CSC_dl_for_check.scala 414:32:@445.4]
  assign _T_1015 = reg2dp_y_extension != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 415:61:@447.4]
  assign _T_1063 = _T_1023 != 7'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 448:37:@484.4]
  assign _T_1064 = ~ _T_1063; // @[NV_NVDLA_CSC_dl_for_check.scala 448:24:@485.4]
  assign _T_1066 = _T_1007 != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 448:56:@486.4]
  assign _T_1067 = ~ _T_1066; // @[NV_NVDLA_CSC_dl_for_check.scala 448:44:@487.4]
  assign _T_1068 = _T_1064 & _T_1067; // @[NV_NVDLA_CSC_dl_for_check.scala 448:42:@488.4]
  assign _T_1070 = _T_996 != 5'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 448:75:@489.4]
  assign _T_1071 = ~ _T_1070; // @[NV_NVDLA_CSC_dl_for_check.scala 448:63:@490.4]
  assign _T_1072 = _T_1068 & _T_1071; // @[NV_NVDLA_CSC_dl_for_check.scala 448:61:@491.4]
  assign _T_1074 = _T_1072 ? 1'h0 : _T_1052; // @[NV_NVDLA_CSC_dl_for_check.scala 448:22:@492.4]
  assign _T_1075 = _T_959 ? 1'h1 : _T_1074; // @[NV_NVDLA_CSC_dl_for_check.scala 447:22:@493.4]
  assign _T_1016 = _T_1015 & _T_1075; // @[NV_NVDLA_CSC_dl_for_check.scala 415:66:@448.4]
  assign _T_1017 = _T_347 | _T_1016; // @[NV_NVDLA_CSC_dl_for_check.scala 415:33:@449.4]
  assign _T_1018 = _T_347 | _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 417:31:@451.6]
  assign _T_1020 = _T_1018 ? 2'h0 : _T_1012; // @[NV_NVDLA_CSC_dl_for_check.scala 417:21:@452.6]
  assign _GEN_65 = _T_1017 ? _T_1020 : _T_1007; // @[NV_NVDLA_CSC_dl_for_check.scala 416:23:@450.4]
  assign _T_1029 = _T_1023 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 425:33:@458.4]
  assign _T_1030 = _T_1023 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 425:33:@459.4]
  assign _T_1031 = _T_1030 == _T_983; // @[NV_NVDLA_CSC_dl_for_check.scala 426:51:@460.4]
  assign _T_1032 = _T_1004 & _T_1031; // @[NV_NVDLA_CSC_dl_for_check.scala 426:33:@461.4]
  assign _T_1033 = _T_1032 & _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 427:34:@463.4]
  assign _T_1034 = _T_1075 & _T_1004; // @[NV_NVDLA_CSC_dl_for_check.scala 428:52:@465.4]
  assign _T_1035 = _T_347 | _T_1034; // @[NV_NVDLA_CSC_dl_for_check.scala 428:34:@466.4]
  assign _T_1037 = ~ _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 432:41:@468.6]
  assign _T_1038 = _T_1032 & _T_1037; // @[NV_NVDLA_CSC_dl_for_check.scala 432:39:@469.6]
  assign _T_1041 = _T_1033 ? 7'h0 : _T_1030; // @[NV_NVDLA_CSC_dl_for_check.scala 433:22:@470.6]
  assign _T_1042 = _T_1038 ? 7'h0 : _T_1041; // @[NV_NVDLA_CSC_dl_for_check.scala 432:22:@471.6]
  assign _T_1043 = _T_347 ? 7'h0 : _T_1042; // @[NV_NVDLA_CSC_dl_for_check.scala 431:22:@472.6]
  assign _GEN_66 = _T_1035 ? _T_1043 : _T_1023; // @[NV_NVDLA_CSC_dl_for_check.scala 430:24:@467.4]
  assign _T_1060 = _T_959 | _T_1046; // @[NV_NVDLA_CSC_dl_for_check.scala 446:27:@482.4]
  assign _T_1055 = _T_1060 & _T_1032; // @[NV_NVDLA_CSC_dl_for_check.scala 443:49:@479.4]
  assign _T_1058 = _T_959 ? 1'h1 : _T_1046; // @[NV_NVDLA_CSC_dl_for_check.scala 444:32:@480.4]
  assign _T_1059 = _T_1055 ? 1'h0 : _T_1058; // @[NV_NVDLA_CSC_dl_for_check.scala 443:33:@481.4]
  assign _T_1080 = {1'h0,_T_982}; // @[Cat.scala 30:58:@499.4]
  assign _GEN_67 = _T_1075 ? _T_1080 : _T_1078; // @[NV_NVDLA_CSC_dl_for_check.scala 458:21:@500.4]
  assign _GEN_683 = {{10'd0}, _T_625}; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@505.4]
  assign _T_1087 = _T_1083 + _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@505.4]
  assign _T_1088 = _T_1083 + _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@506.4]
  assign _T_1089 = _T_1004 & _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 469:29:@507.4]
  assign _T_1090 = _T_1083 >= _T_474; // @[NV_NVDLA_CSC_dl_for_check.scala 469:61:@508.4]
  assign _T_1091 = _T_1089 & _T_1090; // @[NV_NVDLA_CSC_dl_for_check.scala 469:44:@509.4]
  assign _T_1094 = ~ _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 472:43:@512.4]
  assign _T_1095 = _T_1033 & _T_1094; // @[NV_NVDLA_CSC_dl_for_check.scala 472:41:@513.4]
  assign _T_1096 = _T_1091 ? {{9'd0}, _T_365} : _T_1088; // @[NV_NVDLA_CSC_dl_for_check.scala 473:26:@514.4]
  assign _T_1097 = _T_1095 ? _T_1086 : _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 472:26:@515.4]
  assign _T_1098 = _T_347 ? {{9'd0}, _T_365} : _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 471:26:@516.4]
  assign _T_1100 = _T_1034 & _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 474:70:@518.4]
  assign _T_1101 = _T_347 | _T_1100; // @[NV_NVDLA_CSC_dl_for_check.scala 474:37:@519.4]
  assign _T_1102 = _T_1075 & _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 475:55:@520.4]
  assign _T_1103 = _T_1102 & _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 475:71:@521.4]
  assign _T_1104 = _T_347 | _T_1103; // @[NV_NVDLA_CSC_dl_for_check.scala 475:37:@522.4]
  assign _GEN_68 = _T_1101 ? _T_1098 : _T_1083; // @[NV_NVDLA_CSC_dl_for_check.scala 477:27:@523.4]
  assign _GEN_69 = _T_1104 ? _T_1098 : _T_1086; // @[NV_NVDLA_CSC_dl_for_check.scala 480:27:@526.4]
  assign _T_1108 = _T_1107 == _T_583; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@530.4]
  assign _T_1110 = _T_1102 & _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 488:70:@532.4]
  assign _T_1111 = _T_347 | _T_1110; // @[NV_NVDLA_CSC_dl_for_check.scala 488:36:@533.4]
  assign _T_1115 = _T_1107 + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@535.6]
  assign _T_1116 = _T_1107 + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@536.6]
  assign _T_1117 = _T_986 ? 11'h0 : _T_1116; // @[NV_NVDLA_CSC_dl_for_check.scala 492:24:@537.6]
  assign _T_1118 = _T_347 ? 11'h0 : _T_1117; // @[NV_NVDLA_CSC_dl_for_check.scala 491:24:@538.6]
  assign _GEN_70 = _T_1111 ? _T_1118 : _T_1107; // @[NV_NVDLA_CSC_dl_for_check.scala 490:26:@534.4]
  assign _GEN_684 = {{8'd0}, reg2dp_pad_left}; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@550.4]
  assign _T_1147 = 13'h0 - _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@550.4]
  assign _T_1148 = $unsigned(_T_1147); // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@551.4]
  assign _T_1149 = _T_352 ? 14'h0 : _T_1148; // @[NV_NVDLA_CSC_dl_for_check.scala 507:26:@552.4]
  assign _GEN_685 = {{10'd0}, _T_632}; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@553.4]
  assign _T_1150 = _T_1121 + _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@553.4]
  assign _T_1151 = _T_1121 + _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@554.4]
  assign _T_1154 = _T_1091 ? _T_1149 : _T_1151; // @[NV_NVDLA_CSC_dl_for_check.scala 514:25:@557.4]
  assign _T_1155 = _T_1095 ? _T_1124 : _T_1154; // @[NV_NVDLA_CSC_dl_for_check.scala 513:25:@558.4]
  assign _T_1156 = _T_347 ? _T_1149 : _T_1155; // @[NV_NVDLA_CSC_dl_for_check.scala 512:25:@559.4]
  assign _GEN_686 = {{1'd0}, _T_980}; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@560.4]
  assign _T_1157 = _GEN_686 * _T_691; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@560.4]
  assign _GEN_687 = {{3'd0}, _T_1157}; // @[NV_NVDLA_CSC_dl_for_check.scala 517:33:@561.4]
  assign _T_1158 = _T_1121 + _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 517:33:@561.4]
  assign _T_1159 = _T_1121 + _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 517:33:@562.4]
  assign _T_1162 = _T_548[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 518:96:@565.4]
  assign _T_1163 = ~ _T_1162; // @[NV_NVDLA_CSC_dl_for_check.scala 518:86:@566.4]
  assign _T_1164 = _T_1100 & _T_1163; // @[NV_NVDLA_CSC_dl_for_check.scala 518:84:@567.4]
  assign _T_1165 = _T_347 | _T_1164; // @[NV_NVDLA_CSC_dl_for_check.scala 518:36:@568.4]
  assign _T_1168 = _T_548[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 519:99:@571.4]
  assign _T_1169 = ~ _T_1168; // @[NV_NVDLA_CSC_dl_for_check.scala 519:89:@572.4]
  assign _T_1170 = _T_1103 & _T_1169; // @[NV_NVDLA_CSC_dl_for_check.scala 519:87:@573.4]
  assign _T_1171 = _T_347 | _T_1170; // @[NV_NVDLA_CSC_dl_for_check.scala 519:36:@574.4]
  assign _T_1173 = _T_1013 ? _T_670 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 522:26:@575.4]
  assign _T_1176 = _T_387 == 6'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 524:79:@577.4]
  assign _T_1180 = _T_766 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@580.4]
  assign _T_1181 = _T_766 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@581.4]
  assign _T_1182 = _T_1176 ? _T_766 : _T_1181; // @[NV_NVDLA_CSC_dl_for_check.scala 524:27:@582.4]
  assign _T_1183 = _T_986 & _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 526:37:@583.4]
  assign _T_1185 = _T_985 & _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 527:35:@584.4]
  assign _T_1187 = _T_1136 + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 527:66:@585.4]
  assign _T_1188 = _T_1136 + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 527:66:@586.4]
  assign _T_1189 = _T_1185 ? _T_1188 : _T_1136; // @[NV_NVDLA_CSC_dl_for_check.scala 527:22:@587.4]
  assign _T_1190 = _T_1183 ? 13'h2 : _T_1189; // @[NV_NVDLA_CSC_dl_for_check.scala 526:22:@588.4]
  assign _GEN_688 = {{6'd0}, _T_1182}; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@590.4]
  assign _T_1191 = _T_1136 >= _GEN_688; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@590.4]
  assign _T_1192 = _T_1033 & _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 533:39:@591.4]
  assign _T_1193 = _T_1192 & _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 533:54:@592.4]
  assign _T_1194 = _T_1193 & _T_1091; // @[NV_NVDLA_CSC_dl_for_check.scala 533:71:@593.4]
  assign _T_1197 = ~ _T_1091; // @[NV_NVDLA_CSC_dl_for_check.scala 534:73:@596.4]
  assign _T_1198 = _T_1193 & _T_1197; // @[NV_NVDLA_CSC_dl_for_check.scala 534:71:@597.4]
  assign _GEN_689 = {{4'd0}, _T_684}; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@598.4]
  assign _T_1199 = _T_1133 + _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@598.4]
  assign _T_1200 = _T_1133 + _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@599.4]
  assign _T_1202 = _T_1192 & _T_1191; // @[NV_NVDLA_CSC_dl_for_check.scala 535:54:@601.4]
  assign _GEN_690 = {{9'd0}, _T_663}; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@602.4]
  assign _T_1203 = _T_1130 + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@602.4]
  assign _T_1204 = _T_1130 + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@603.4]
  assign _T_1206 = ~ _T_1191; // @[NV_NVDLA_CSC_dl_for_check.scala 536:56:@605.4]
  assign _T_1207 = _T_1192 & _T_1206; // @[NV_NVDLA_CSC_dl_for_check.scala 536:54:@606.4]
  assign _T_1209 = _T_1130 + 16'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 536:91:@607.4]
  assign _T_1210 = _T_1130 + 16'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 536:91:@608.4]
  assign _T_1211 = ~ _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 537:41:@609.4]
  assign _T_1212 = _T_1033 & _T_1211; // @[NV_NVDLA_CSC_dl_for_check.scala 537:39:@610.4]
  assign _GEN_691 = {{8'd0}, _T_1173}; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@611.4]
  assign _T_1213 = _T_1127 + _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@611.4]
  assign _T_1214 = _T_1127 + _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@612.4]
  assign _T_1215 = _T_1212 ? _T_1130 : _T_1214; // @[NV_NVDLA_CSC_dl_for_check.scala 537:24:@613.4]
  assign _T_1216 = _T_1207 ? _T_1210 : _T_1215; // @[NV_NVDLA_CSC_dl_for_check.scala 536:24:@614.4]
  assign _T_1217 = _T_1202 ? _T_1204 : _T_1216; // @[NV_NVDLA_CSC_dl_for_check.scala 535:24:@615.4]
  assign _T_1218 = _T_1198 ? _T_1200 : _T_1217; // @[NV_NVDLA_CSC_dl_for_check.scala 534:24:@616.4]
  assign _T_1219 = _T_1194 ? {{9'd0}, _T_656} : _T_1218; // @[NV_NVDLA_CSC_dl_for_check.scala 533:24:@617.4]
  assign _T_1220 = _T_432 ? {{9'd0}, _T_656} : _T_1219; // @[NV_NVDLA_CSC_dl_for_check.scala 532:24:@618.4]
  assign _T_1226 = _T_1127[15:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 539:68:@620.4]
  assign _T_1227 = {5'h0,_T_1226}; // @[Cat.scala 30:58:@621.4]
  assign _T_1238 = _T_548[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 542:68:@632.4]
  assign _T_1239 = _T_1075 & _T_1238; // @[NV_NVDLA_CSC_dl_for_check.scala 542:57:@633.4]
  assign _T_1240 = _T_1239 & _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 542:72:@634.4]
  assign _T_1241 = _T_1240 & _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 542:88:@635.4]
  assign _T_1242 = _T_1241 & _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 542:103:@636.4]
  assign _T_1243 = _T_432 | _T_1242; // @[NV_NVDLA_CSC_dl_for_check.scala 542:39:@637.4]
  assign _T_1245 = _T_1162 & _T_959; // @[NV_NVDLA_CSC_dl_for_check.scala 544:42:@639.4]
  assign _T_1248 = _T_1141 ? 1'h0 : _T_1144; // @[NV_NVDLA_CSC_dl_for_check.scala 544:74:@640.4]
  assign _T_1249 = _T_1245 ? 1'h1 : _T_1248; // @[NV_NVDLA_CSC_dl_for_check.scala 544:28:@641.4]
  assign _T_1251 = _T_1162 & _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 545:36:@643.4]
  assign _T_1252 = _T_1249 | _T_1144; // @[NV_NVDLA_CSC_dl_for_check.scala 545:72:@644.4]
  assign _T_1253 = _T_1251 & _T_1252; // @[NV_NVDLA_CSC_dl_for_check.scala 545:51:@645.4]
  assign _GEN_71 = _T_1165 ? _T_1156 : _T_1121; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@646.4]
  assign _GEN_72 = _T_1165 ? _T_1220 : _T_1127; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@646.4]
  assign _GEN_73 = _T_1171 ? _T_1156 : _T_1124; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@650.4]
  assign _GEN_74 = _T_1171 ? _T_1220 : _T_1130; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@650.4]
  assign _GEN_75 = _T_1243 ? _T_1220 : _T_1133; // @[NV_NVDLA_CSC_dl_for_check.scala 555:26:@654.4]
  assign _GEN_692 = {{9'd0}, reg2dp_pad_top}; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@659.4]
  assign _T_1261 = 14'h0 - _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@659.4]
  assign _T_1262 = $unsigned(_T_1261); // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@660.4]
  assign _T_1263 = _T_1262[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@661.4]
  assign _GEN_693 = {{10'd0}, _T_639}; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@662.4]
  assign _T_1264 = _T_1256 + _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@662.4]
  assign _T_1265 = _T_1256 + _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@663.4]
  assign _T_1266 = _T_1033 & _T_987; // @[NV_NVDLA_CSC_dl_for_check.scala 566:52:@664.4]
  assign _T_1267 = _T_347 | _T_1266; // @[NV_NVDLA_CSC_dl_for_check.scala 566:35:@665.4]
  assign _T_1270 = _T_1091 ? _T_1265 : _T_1256; // @[NV_NVDLA_CSC_dl_for_check.scala 568:25:@668.4]
  assign _T_1271 = _T_1095 ? _T_1259 : _T_1270; // @[NV_NVDLA_CSC_dl_for_check.scala 567:25:@669.4]
  assign _T_1272 = _T_1267 ? _T_1263 : _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 566:25:@670.4]
  assign _T_1275 = _T_1095 | _T_1091; // @[NV_NVDLA_CSC_dl_for_check.scala 569:91:@673.4]
  assign _T_1276 = _T_1075 & _T_1275; // @[NV_NVDLA_CSC_dl_for_check.scala 569:54:@674.4]
  assign _T_1277 = _T_347 | _T_1276; // @[NV_NVDLA_CSC_dl_for_check.scala 569:36:@675.4]
  assign _GEN_694 = {{1'd0}, _T_981}; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@679.4]
  assign _T_1281 = _GEN_694 * _T_698; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@679.4]
  assign _GEN_695 = {{3'd0}, _T_1281}; // @[NV_NVDLA_CSC_dl_for_check.scala 572:33:@680.4]
  assign _T_1282 = _T_1256 + _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 572:33:@680.4]
  assign _T_1283 = _T_1256 + _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 572:33:@681.4]
  assign _GEN_696 = {{12'd0}, _T_1007}; // @[NV_NVDLA_CSC_dl_for_check.scala 572:51:@682.4]
  assign _T_1284 = _T_1283 + _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 572:51:@682.4]
  assign _T_1285 = _T_1283 + _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 572:51:@683.4]
  assign _GEN_76 = _T_1277 ? _T_1272 : _T_1256; // @[NV_NVDLA_CSC_dl_for_check.scala 574:26:@684.4]
  assign _GEN_77 = _T_1104 ? _T_1272 : _T_1259; // @[NV_NVDLA_CSC_dl_for_check.scala 575:26:@687.4]
  assign _T_1286 = _T_1159[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 578:39:@690.4]
  assign _GEN_697 = {{1'd0}, _T_569}; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@691.4]
  assign _T_1287 = _T_1159 > _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@691.4]
  assign _T_1288 = _T_1286 | _T_1287; // @[NV_NVDLA_CSC_dl_for_check.scala 578:44:@692.4]
  assign _T_1289 = _T_1285[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 578:92:@693.4]
  assign _T_1290 = _T_1288 | _T_1289; // @[NV_NVDLA_CSC_dl_for_check.scala 578:78:@694.4]
  assign _GEN_698 = {{1'd0}, _T_576}; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@695.4]
  assign _T_1291 = _T_1285 > _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@695.4]
  assign _T_1292 = _T_1290 | _T_1291; // @[NV_NVDLA_CSC_dl_for_check.scala 578:97:@696.4]
  assign _T_1305 = _T_1289 | _T_1291; // @[NV_NVDLA_CSC_dl_for_check.scala 581:42:@706.4]
  assign _T_1415 = _T_548[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 666:33:@792.4]
  assign _T_1416 = ~ _T_1108; // @[NV_NVDLA_CSC_dl_for_check.scala 667:24:@793.4]
  assign _T_1418 = _T_1159[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 667:77:@794.4]
  assign _T_1419 = {2'h0,_T_1418}; // @[Cat.scala 30:58:@795.4]
  assign _T_1421 = _T_1080 > 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 668:38:@796.4]
  assign _T_1426 = _T_1159[12:1]; // @[NV_NVDLA_CSC_dl_for_check.scala 669:54:@799.4]
  assign _T_1427 = {3'h0,_T_1426}; // @[Cat.scala 30:58:@800.4]
  assign _T_1428 = _T_1421 ? _T_1419 : _T_1427; // @[NV_NVDLA_CSC_dl_for_check.scala 668:23:@801.4]
  assign _T_1429 = _T_1416 ? _T_1419 : _T_1428; // @[NV_NVDLA_CSC_dl_for_check.scala 667:23:@802.4]
  assign _T_1430 = _T_1415 ? _T_1227 : _T_1429; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@803.4]
  assign _T_1431 = _T_1430[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 678:24:@805.4]
  assign _T_1308 = _T_1431[13:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 585:32:@708.4]
  assign _GEN_700 = {{3'd0}, _T_1308}; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@709.4]
  assign _T_1309 = _GEN_700 > _T_712; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@709.4]
  assign _T_1310 = _T_548[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 586:34:@710.4]
  assign _T_1311 = _T_1310 ? _T_1305 : _T_1292; // @[NV_NVDLA_CSC_dl_for_check.scala 586:24:@711.4]
  assign _T_1312 = _T_548[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 587:29:@712.4]
  assign _T_1313 = _T_1312 & _T_1309; // @[NV_NVDLA_CSC_dl_for_check.scala 587:33:@713.4]
  assign _T_1314 = ~ _T_1311; // @[NV_NVDLA_CSC_dl_for_check.scala 588:39:@714.4]
  assign _T_1315 = _T_1075 & _T_1314; // @[NV_NVDLA_CSC_dl_for_check.scala 588:37:@715.4]
  assign _T_1316 = ~ _T_1313; // @[NV_NVDLA_CSC_dl_for_check.scala 588:56:@716.4]
  assign _T_1317 = _T_1315 & _T_1316; // @[NV_NVDLA_CSC_dl_for_check.scala 588:54:@717.4]
  assign _T_1318 = _T_548[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 591:37:@718.4]
  assign _T_1319 = ~ _T_1318; // @[NV_NVDLA_CSC_dl_for_check.scala 591:27:@719.4]
  assign _T_1320 = _T_1107[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 591:54:@720.4]
  assign _T_1321 = _T_1319 ? _T_1320 : _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 591:26:@721.4]
  assign _T_1322 = _T_1159[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 592:35:@722.4]
  assign _T_1324 = _T_1007 == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 593:55:@723.4]
  assign _T_1325 = _T_1075 & _T_1324; // @[NV_NVDLA_CSC_dl_for_check.scala 593:42:@724.4]
  assign _T_1326 = _T_1032 & _T_1060; // @[NV_NVDLA_CSC_dl_for_check.scala 596:42:@726.4]
  assign _T_1330 = {_T_988,_T_986,_T_1326,_T_959,_T_996}; // @[Cat.scala 30:58:@730.4]
  assign _T_1361 = _T_989 & _T_1032; // @[NV_NVDLA_CSC_dl_for_check.scala 623:38:@750.6]
  assign _T_1362 = _T_1361 & _T_1060; // @[NV_NVDLA_CSC_dl_for_check.scala 623:56:@751.6]
  assign _GEN_78 = _T_1075 ? _T_1322 : _T_1336; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_79 = _T_1075 ? _T_1007 : _T_1339; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_80 = _T_1075 ? _T_1321 : _T_1342; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_81 = _T_1075 ? _T_1108 : _T_1345; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_82 = _T_1075 ? _T_1075 : _T_1348; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_83 = _T_1075 ? _T_984 : _T_1351; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_84 = _T_1075 ? _T_1330 : _T_1357; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_85 = _T_1075 ? _T_1362 : _T_1360; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_86 = _T_1075 ? _T_1249 : _T_1144; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_87 = _T_1075 ? _T_1253 : _T_1141; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@742.4]
  assign _GEN_88 = _T_1325 ? _T_959 : _T_1354; // @[NV_NVDLA_CSC_dl_for_check.scala 627:26:@756.4]
  assign _T_1384 = _T_548[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 644:32:@766.4]
  assign _T_1385 = ~ _T_1384; // @[NV_NVDLA_CSC_dl_for_check.scala 644:22:@767.4]
  assign _T_1386 = _T_562[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 644:49:@768.4]
  assign _T_1388 = _T_1385 ? _T_1386 : 12'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 644:21:@769.4]
  assign _T_1390 = _T_1033 & _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 646:34:@770.4]
  assign _GEN_701 = {{1'd0}, _T_1388}; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@771.4]
  assign _T_1392 = _T_1365 + _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@771.4]
  assign _T_1393 = _T_1365 + _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@772.4]
  assign _T_1394 = _T_1390 ? 13'h0 : _T_1393; // @[NV_NVDLA_CSC_dl_for_check.scala 646:19:@773.4]
  assign _T_1395 = _T_347 ? 13'h0 : _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 645:19:@774.4]
  assign _T_1399 = _T_1365 != _T_1368; // @[NV_NVDLA_CSC_dl_for_check.scala 648:31:@778.4]
  assign _GEN_702 = {{2'd0}, _T_495}; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@779.4]
  assign _T_1400 = _T_1256 * _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@779.4]
  assign _T_1401 = _T_1400[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 651:50:@780.4]
  assign _GEN_703 = {{7'd0}, _T_981}; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@781.4]
  assign _T_1402 = _GEN_703 * _T_502; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@781.4]
  assign _T_1403 = _T_1402[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 652:49:@782.4]
  assign _GEN_704 = {{10'd0}, _T_996}; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@783.4]
  assign _T_1404 = _GEN_704 * _T_719; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@783.4]
  assign _T_1405 = _T_1404[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 653:47:@784.4]
  assign _GEN_705 = {{13'd0}, _T_1007}; // @[NV_NVDLA_CSC_dl_for_check.scala 654:47:@785.4]
  assign _T_1407 = _GEN_705 * _T_726; // @[NV_NVDLA_CSC_dl_for_check.scala 654:47:@785.4]
  assign _T_1408 = _T_347 ? 17'h0 : _T_1407; // @[NV_NVDLA_CSC_dl_for_check.scala 654:21:@786.4]
  assign _T_1409 = _T_1408[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 654:65:@787.4]
  assign _T_1410 = _T_548[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 655:45:@788.4]
  assign _T_1411 = _T_347 | _T_1410; // @[NV_NVDLA_CSC_dl_for_check.scala 655:34:@789.4]
  assign _T_1412 = {_T_1411,_T_1075}; // @[Cat.scala 30:58:@790.4]
  assign _GEN_89 = _T_1111 ? _T_1395 : _T_1365; // @[NV_NVDLA_CSC_dl_for_check.scala 682:20:@807.4]
  assign _GEN_90 = _T_1399 ? _T_1365 : _T_1368; // @[NV_NVDLA_CSC_dl_for_check.scala 685:23:@810.4]
  assign _T_1432 = _T_1412[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 688:19:@813.4]
  assign _GEN_91 = _T_1432 ? _T_1401 : _T_1371; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@814.4]
  assign _GEN_92 = _T_1432 ? _T_1403 : _T_1374; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@814.4]
  assign _GEN_93 = _T_1432 ? _T_1405 : _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@814.4]
  assign _T_1433 = _T_1412[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 693:19:@819.4]
  assign _GEN_94 = _T_1433 ? _T_1409 : _T_1380; // @[NV_NVDLA_CSC_dl_for_check.scala 693:23:@820.4]
  assign _GEN_95 = _T_1075 ? _T_1431 : {{1'd0}, _T_1383}; // @[NV_NVDLA_CSC_dl_for_check.scala 696:20:@823.4]
  assign _T_1539 = _T_1371 + _T_1374; // @[NV_NVDLA_CSC_dl_for_check.scala 720:29:@851.4]
  assign _T_1540 = _T_1371 + _T_1374; // @[NV_NVDLA_CSC_dl_for_check.scala 720:29:@852.4]
  assign _T_1541 = _T_1540 + _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 720:43:@853.4]
  assign _T_1542 = _T_1540 + _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 720:43:@854.4]
  assign _T_1543 = _T_1542 + _T_1380; // @[NV_NVDLA_CSC_dl_for_check.scala 720:57:@855.4]
  assign _T_1544 = _T_1542 + _T_1380; // @[NV_NVDLA_CSC_dl_for_check.scala 720:57:@856.4]
  assign _GEN_706 = {{2'd0}, _T_1368}; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@857.4]
  assign _T_1545 = _T_793 + _GEN_706; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@857.4]
  assign _T_1546 = _T_793 + _GEN_706; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@858.4]
  assign _GEN_707 = {{2'd0}, _T_1544}; // @[NV_NVDLA_CSC_dl_for_check.scala 721:52:@859.4]
  assign _T_1547 = _T_1546 + _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 721:52:@859.4]
  assign _T_1548 = _T_1546 + _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 721:52:@860.4]
  assign _GEN_708 = {{2'd0}, _T_1383}; // @[NV_NVDLA_CSC_dl_for_check.scala 721:64:@861.4]
  assign _T_1549 = _T_1548 + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 721:64:@861.4]
  assign _T_1550 = _T_1548 + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 721:64:@862.4]
  assign _T_1557 = _T_1550 >= _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 722:45:@865.4]
  assign _T_1564 = _T_1550 - _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@868.4]
  assign _T_1565 = $unsigned(_T_1564); // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@869.4]
  assign _T_1566 = _T_1565[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@870.4]
  assign _T_1567 = _T_347 | _T_1348; // @[NV_NVDLA_CSC_dl_for_check.scala 724:35:@871.4]
  assign _T_1573 = _T_1557 ? _T_1566 : _T_1550; // @[NV_NVDLA_CSC_dl_for_check.scala 725:25:@873.4]
  assign _T_1574 = _T_1567 ? 15'h1fff : _T_1573; // @[NV_NVDLA_CSC_dl_for_check.scala 724:25:@874.4]
  assign _T_1598 = 2'h3 == _T_1339; // @[Mux.scala 46:19:@884.4]
  assign _T_1599 = _T_1598 ? _T_1476_3 : 13'h0; // @[Mux.scala 46:16:@885.4]
  assign _T_1600 = 2'h2 == _T_1339; // @[Mux.scala 46:19:@886.4]
  assign _T_1601 = _T_1600 ? _T_1476_2 : _T_1599; // @[Mux.scala 46:16:@887.4]
  assign _T_1602 = 2'h1 == _T_1339; // @[Mux.scala 46:19:@888.4]
  assign _T_1603 = _T_1602 ? _T_1476_1 : _T_1601; // @[Mux.scala 46:16:@889.4]
  assign _T_1604 = 2'h0 == _T_1339; // @[Mux.scala 46:19:@890.4]
  assign _T_1605 = _T_1604 ? _T_1476_0 : _T_1603; // @[Mux.scala 46:16:@891.4]
  assign _GEN_712 = {{2'd0}, _T_1605}; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@892.4]
  assign _T_1606 = _GEN_712 != _T_1574; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@892.4]
  assign _T_1607 = _T_1606 | _T_1144; // @[NV_NVDLA_CSC_dl_for_check.scala 732:85:@893.4]
  assign _T_1608 = _T_1333 & _T_1607; // @[NV_NVDLA_CSC_dl_for_check.scala 732:43:@894.4]
  assign _T_1609 = _T_1333 | _T_1348; // @[NV_NVDLA_CSC_dl_for_check.scala 734:38:@895.4]
  assign _T_1611 = _T_1339 == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@896.4]
  assign _T_1612 = _T_1609 & _T_1611; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@897.4]
  assign _T_1613 = _T_347 | _T_1612; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@898.4]
  assign _T_1616 = _T_1339 == 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@900.4]
  assign _T_1617 = _T_1609 & _T_1616; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@901.4]
  assign _T_1618 = _T_347 | _T_1617; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@902.4]
  assign _T_1621 = _T_1339 == 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@904.4]
  assign _T_1622 = _T_1609 & _T_1621; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@905.4]
  assign _T_1623 = _T_347 | _T_1622; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@906.4]
  assign _T_1626 = _T_1339 == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@908.4]
  assign _T_1627 = _T_1609 & _T_1626; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@909.4]
  assign _T_1628 = _T_347 | _T_1627; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@910.4]
  assign _GEN_96 = _T_1613 ? _T_1574 : {{2'd0}, _T_1476_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@916.4]
  assign _GEN_97 = _T_1618 ? _T_1574 : {{2'd0}, _T_1476_1}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@919.4]
  assign _GEN_98 = _T_1623 ? _T_1574 : {{2'd0}, _T_1476_2}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@922.4]
  assign _GEN_99 = _T_1628 ? _T_1574 : {{2'd0}, _T_1476_3}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@925.4]
  assign _T_1639 = _T_347 | _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 747:14:@929.4]
  assign _GEN_100 = _T_1639 ? _T_1574 : _T_1502; // @[NV_NVDLA_CSC_dl_for_check.scala 747:34:@930.4]
  assign _GEN_101 = _T_1052 ? _T_1336 : _T_1511; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_102 = _T_1052 ? _T_1339 : _T_1514; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_103 = _T_1052 ? _T_1342 : _T_1517; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_104 = _T_1052 ? _T_1345 : _T_1520; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_105 = _T_1052 ? _T_1078 : _T_1523; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_106 = _T_1052 ? _T_1348 : _T_1526; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_107 = _T_1052 ? _T_1351 : _T_1529; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_108 = _T_1052 ? _T_1354 : _T_1532; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_109 = _T_1052 ? _T_1360 : _T_1535; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _GEN_110 = _T_1052 ? _T_1357 : {{8'd0}, _T_1052}; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@937.4]
  assign _T_1649 = {1'h0,_T_1520,_T_1517,_T_1514,_T_1511}; // @[Cat.scala 30:58:@957.4]
  assign _T_1655 = {_T_1538,_T_1535,_T_1532,_T_1526,_T_1529,_T_1523,_T_1649}; // @[Cat.scala 30:58:@963.4]
  assign _GEN_111 = _T_1505 ? _T_1655 : _T_1680; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1005.4]
  assign _GEN_114 = _T_1660 ? _T_1680 : _T_1683; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1014.4]
  assign _GEN_117 = _T_1663 ? _T_1683 : _T_1686; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1023.4]
  assign _GEN_120 = _T_1666 ? _T_1686 : _T_1689; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1032.4]
  assign _GEN_123 = _T_1669 ? _T_1689 : _T_1692; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1041.4]
  assign _GEN_126 = _T_1672 ? _T_1692 : _T_1695; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1050.4]
  assign _T_1756 = _T_1695[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 816:41:@1058.4]
  assign _T_1757 = _T_1695[3:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 817:41:@1059.4]
  assign _T_1758 = _T_1695[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 818:41:@1060.4]
  assign _T_1759 = _T_1695[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 819:42:@1061.4]
  assign _T_1760 = _T_1695[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 820:41:@1062.4]
  assign _T_1761 = _T_1695[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 821:45:@1063.4]
  assign _T_1764 = _T_1695[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 824:39:@1066.4]
  assign _T_1765 = _T_1695[28:20]; // @[NV_NVDLA_CSC_dl_for_check.scala 825:40:@1067.4]
  assign _T_1822 = _T_548[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 855:69:@1095.4]
  assign _T_1823 = _T_1822 & sc2buf_dat_rd_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 855:74:@1096.4]
  assign _T_1824 = ~ _T_1768; // @[NV_NVDLA_CSC_dl_for_check.scala 855:90:@1097.4]
  assign _T_1825 = _T_1823 & _T_1824; // @[NV_NVDLA_CSC_dl_for_check.scala 855:88:@1098.4]
  assign _T_1865 = sc2buf_dat_rd_valid ? 1'h0 : _T_1768; // @[NV_NVDLA_CSC_dl_for_check.scala 870:22:@1132.4]
  assign _T_1879 = sc2buf_dat_rd_valid ? _T_1768 : _T_1780; // @[NV_NVDLA_CSC_dl_for_check.scala 874:48:@1143.4]
  assign _T_1880 = _T_1825 ? 1'h0 : _T_1879; // @[NV_NVDLA_CSC_dl_for_check.scala 874:22:@1144.4]
  assign _T_1957 = {_T_1765,_T_1764,_T_1761,_T_1760,1'h0,_T_1759,_T_1758,_T_1757,_T_1756}; // @[Cat.scala 30:58:@1211.4]
  assign _GEN_137 = _T_1675 ? _T_1957 : _T_1939; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1214.4]
  assign _GEN_138 = _T_1925 ? _T_1939 : _T_1942; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1218.4]
  assign _GEN_139 = _T_1928 ? _T_1942 : _T_1945; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1222.4]
  assign _GEN_140 = _T_1931 ? _T_1945 : _T_1948; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1226.4]
  assign _T_1986 = _T_1939[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 931:39:@1252.4]
  assign _T_1987 = _T_1942[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 932:39:@1253.4]
  assign _T_1988 = _T_1945[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 933:39:@1254.4]
  assign _T_1989 = _T_1948[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 934:39:@1255.4]
  assign _T_1990 = _T_1939[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 936:38:@1256.4]
  assign _T_1991 = _T_1942[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 937:38:@1257.4]
  assign _T_1992 = _T_1945[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 938:38:@1258.4]
  assign _T_1993 = _T_1948[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 939:38:@1259.4]
  assign _T_1994 = _T_1990[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 941:44:@1260.4]
  assign _T_1995 = _T_1991[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 942:44:@1261.4]
  assign _T_1996 = _T_1992[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 943:44:@1262.4]
  assign _T_1997 = _T_1993[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 944:44:@1263.4]
  assign _T_1998 = _T_1985[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 947:31:@1264.4]
  assign _T_2002 = _T_1985[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 951:31:@1268.4]
  assign _T_2003 = _T_1985[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 952:35:@1269.4]
  assign _T_2013 = sc2buf_dat_rd_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 963:29:@1278.4]
  assign _T_2024 = _T_677 > 7'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 968:50:@1282.4]
  assign _GEN_713 = {{1'd0}, _T_677}; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1283.4]
  assign _T_2026 = _T_1899 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1283.4]
  assign _T_2027 = _T_1899 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1284.4]
  assign _T_2028 = _T_2027 - _T_2013; // @[NV_NVDLA_CSC_dl_for_check.scala 968:133:@1285.4]
  assign _T_2029 = $unsigned(_T_2028); // @[NV_NVDLA_CSC_dl_for_check.scala 968:133:@1286.4]
  assign _T_2030 = _T_2029[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 968:133:@1287.4]
  assign _T_2031 = _T_2024 ? 8'h40 : _T_2030; // @[NV_NVDLA_CSC_dl_for_check.scala 968:29:@1288.4]
  assign _T_2035 = _T_1902 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 969:111:@1290.4]
  assign _T_2036 = _T_1902 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 969:111:@1291.4]
  assign _T_2037 = _T_2036 - 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 969:133:@1292.4]
  assign _T_2038 = $unsigned(_T_2037); // @[NV_NVDLA_CSC_dl_for_check.scala 969:133:@1293.4]
  assign _T_2039 = _T_2038[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 969:133:@1294.4]
  assign _T_2040 = _T_2024 ? 8'h40 : _T_2039; // @[NV_NVDLA_CSC_dl_for_check.scala 969:29:@1295.4]
  assign _T_2044 = _T_1905 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 970:111:@1297.4]
  assign _T_2045 = _T_1905 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 970:111:@1298.4]
  assign _T_2046 = _T_2045 - 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 970:133:@1299.4]
  assign _T_2047 = $unsigned(_T_2046); // @[NV_NVDLA_CSC_dl_for_check.scala 970:133:@1300.4]
  assign _T_2048 = _T_2047[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 970:133:@1301.4]
  assign _T_2049 = _T_2024 ? 8'h40 : _T_2048; // @[NV_NVDLA_CSC_dl_for_check.scala 970:29:@1302.4]
  assign _T_2053 = _T_1908 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 971:111:@1304.4]
  assign _T_2054 = _T_1908 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 971:111:@1305.4]
  assign _T_2055 = _T_2054 - 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 971:133:@1306.4]
  assign _T_2056 = $unsigned(_T_2055); // @[NV_NVDLA_CSC_dl_for_check.scala 971:133:@1307.4]
  assign _T_2057 = _T_2056[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 971:133:@1308.4]
  assign _T_2058 = _T_2024 ? 8'h40 : _T_2057; // @[NV_NVDLA_CSC_dl_for_check.scala 971:29:@1309.4]
  assign _T_2060 = ~ _T_1986; // @[NV_NVDLA_CSC_dl_for_check.scala 980:52:@1310.4]
  assign _T_2061 = _T_1994 & _T_2060; // @[NV_NVDLA_CSC_dl_for_check.scala 980:50:@1311.4]
  assign _T_2062 = _T_1994 & _T_1986; // @[NV_NVDLA_CSC_dl_for_check.scala 981:50:@1312.4]
  assign _T_2067 = _T_2062 ? 8'h40 : _T_2031; // @[NV_NVDLA_CSC_dl_for_check.scala 981:27:@1315.4]
  assign _T_2068 = _T_2061 ? _T_1911 : _T_2067; // @[NV_NVDLA_CSC_dl_for_check.scala 980:27:@1316.4]
  assign _T_2069 = _T_347 ? 8'h40 : _T_2068; // @[NV_NVDLA_CSC_dl_for_check.scala 979:27:@1317.4]
  assign _T_2071 = ~ _T_1987; // @[NV_NVDLA_CSC_dl_for_check.scala 985:52:@1318.4]
  assign _T_2072 = _T_1995 & _T_2071; // @[NV_NVDLA_CSC_dl_for_check.scala 985:50:@1319.4]
  assign _T_2073 = _T_1995 & _T_1987; // @[NV_NVDLA_CSC_dl_for_check.scala 986:50:@1320.4]
  assign _T_2078 = _T_2073 ? 8'h40 : _T_2040; // @[NV_NVDLA_CSC_dl_for_check.scala 986:27:@1323.4]
  assign _T_2079 = _T_2072 ? _T_1914 : _T_2078; // @[NV_NVDLA_CSC_dl_for_check.scala 985:27:@1324.4]
  assign _T_2080 = _T_347 ? 8'h40 : _T_2079; // @[NV_NVDLA_CSC_dl_for_check.scala 984:27:@1325.4]
  assign _T_2082 = ~ _T_1988; // @[NV_NVDLA_CSC_dl_for_check.scala 990:52:@1326.4]
  assign _T_2083 = _T_1996 & _T_2082; // @[NV_NVDLA_CSC_dl_for_check.scala 990:50:@1327.4]
  assign _T_2084 = _T_1996 & _T_1988; // @[NV_NVDLA_CSC_dl_for_check.scala 991:50:@1328.4]
  assign _T_2089 = _T_2084 ? 8'h40 : _T_2049; // @[NV_NVDLA_CSC_dl_for_check.scala 991:27:@1331.4]
  assign _T_2090 = _T_2083 ? _T_1917 : _T_2089; // @[NV_NVDLA_CSC_dl_for_check.scala 990:27:@1332.4]
  assign _T_2091 = _T_347 ? 8'h40 : _T_2090; // @[NV_NVDLA_CSC_dl_for_check.scala 989:27:@1333.4]
  assign _T_2093 = ~ _T_1989; // @[NV_NVDLA_CSC_dl_for_check.scala 995:52:@1334.4]
  assign _T_2094 = _T_1997 & _T_2093; // @[NV_NVDLA_CSC_dl_for_check.scala 995:50:@1335.4]
  assign _T_2095 = _T_1997 & _T_1989; // @[NV_NVDLA_CSC_dl_for_check.scala 996:50:@1336.4]
  assign _T_2100 = _T_2095 ? 8'h40 : _T_2058; // @[NV_NVDLA_CSC_dl_for_check.scala 996:27:@1339.4]
  assign _T_2101 = _T_2094 ? _T_1920 : _T_2100; // @[NV_NVDLA_CSC_dl_for_check.scala 995:27:@1340.4]
  assign _T_2102 = _T_347 ? 8'h40 : _T_2101; // @[NV_NVDLA_CSC_dl_for_check.scala 994:27:@1341.4]
  assign _T_2103 = _T_548[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:46:@1342.4]
  assign _T_2104 = _T_2103 & _T_1925; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:51:@1343.4]
  assign _T_2105 = _T_347 | _T_2104; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:34:@1344.4]
  assign _T_2106 = _T_548[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:46:@1345.4]
  assign _T_2107 = _T_2106 & _T_1928; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:51:@1346.4]
  assign _T_2109 = _T_601 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:87:@1347.4]
  assign _T_2110 = _T_2107 & _T_2109; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:69:@1348.4]
  assign _T_2111 = _T_347 | _T_2110; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:34:@1349.4]
  assign _T_2112 = _T_548[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:46:@1350.4]
  assign _T_2113 = _T_2112 & _T_1931; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:51:@1351.4]
  assign _T_2115 = _T_601 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:87:@1352.4]
  assign _T_2116 = _T_2113 & _T_2115; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:69:@1353.4]
  assign _T_2117 = _T_347 | _T_2116; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:34:@1354.4]
  assign _T_2118 = _T_548[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:46:@1355.4]
  assign _T_2119 = _T_2118 & _T_1934; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:51:@1356.4]
  assign _T_2122 = _T_2119 & _T_2115; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:69:@1358.4]
  assign _T_2123 = _T_347 | _T_2122; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:34:@1359.4]
  assign _T_2124 = _T_548[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:50:@1360.4]
  assign _T_2125 = _T_2124 & _T_1925; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:55:@1361.4]
  assign _T_2126 = _T_2125 & _T_1994; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:73:@1362.4]
  assign _T_2127 = _T_2126 & _T_1986; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:97:@1363.4]
  assign _T_2128 = _T_347 | _T_2127; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:38:@1364.4]
  assign _T_2129 = _T_548[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:50:@1365.4]
  assign _T_2130 = _T_2129 & _T_1928; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:55:@1366.4]
  assign _T_2131 = _T_2130 & _T_1995; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:73:@1367.4]
  assign _T_2132 = _T_2131 & _T_1987; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:97:@1368.4]
  assign _T_2134 = _T_604 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:138:@1369.4]
  assign _T_2135 = _T_2132 & _T_2134; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:120:@1370.4]
  assign _T_2136 = _T_347 | _T_2135; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:38:@1371.4]
  assign _T_2137 = _T_548[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:50:@1372.4]
  assign _T_2138 = _T_2137 & _T_1931; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:55:@1373.4]
  assign _T_2139 = _T_2138 & _T_1996; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:73:@1374.4]
  assign _T_2140 = _T_2139 & _T_1988; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:97:@1375.4]
  assign _T_2142 = _T_604 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:138:@1376.4]
  assign _T_2143 = _T_2140 & _T_2142; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:120:@1377.4]
  assign _T_2144 = _T_347 | _T_2143; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:38:@1378.4]
  assign _T_2145 = _T_548[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:50:@1379.4]
  assign _T_2146 = _T_2145 & _T_1934; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:55:@1380.4]
  assign _T_2147 = _T_2146 & _T_1997; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:73:@1381.4]
  assign _T_2148 = _T_2147 & _T_1989; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:97:@1382.4]
  assign _T_2151 = _T_2148 & _T_2142; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:120:@1384.4]
  assign _T_2152 = _T_347 | _T_2151; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:38:@1385.4]
  assign _GEN_141 = _T_2105 ? _T_2069 : _T_1899; // @[NV_NVDLA_CSC_dl_for_check.scala 1010:24:@1386.4]
  assign _GEN_142 = _T_2111 ? _T_2080 : _T_1902; // @[NV_NVDLA_CSC_dl_for_check.scala 1011:24:@1389.4]
  assign _GEN_143 = _T_2117 ? _T_2091 : _T_1905; // @[NV_NVDLA_CSC_dl_for_check.scala 1012:24:@1392.4]
  assign _GEN_144 = _T_2123 ? _T_2102 : _T_1908; // @[NV_NVDLA_CSC_dl_for_check.scala 1013:24:@1395.4]
  assign _GEN_145 = _T_2128 ? _T_2069 : _T_1911; // @[NV_NVDLA_CSC_dl_for_check.scala 1014:28:@1398.4]
  assign _GEN_146 = _T_2136 ? _T_2080 : _T_1914; // @[NV_NVDLA_CSC_dl_for_check.scala 1015:28:@1401.4]
  assign _GEN_147 = _T_2144 ? _T_2091 : _T_1917; // @[NV_NVDLA_CSC_dl_for_check.scala 1016:28:@1404.4]
  assign _GEN_148 = _T_2152 ? _T_2102 : _T_1920; // @[NV_NVDLA_CSC_dl_for_check.scala 1017:28:@1407.4]
  assign _T_2153 = _T_705[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:55:@1410.4]
  assign _T_2156 = {_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153}; // @[Cat.scala 30:58:@1413.4]
  assign _T_2157 = {_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2156}; // @[Cat.scala 30:58:@1414.4]
  assign _T_2158 = {_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2153,_T_2156,_T_2157}; // @[Cat.scala 30:58:@1415.4]
  assign _T_2159 = {_T_2158,_T_2158}; // @[Cat.scala 30:58:@1416.4]
  assign _T_2160 = _T_1768 ? _T_2159 : _T_1791; // @[NV_NVDLA_CSC_dl_for_check.scala 1028:23:@1417.4]
  assign _T_2164 = _T_1780 ? _T_2159 : _T_1799; // @[NV_NVDLA_CSC_dl_for_check.scala 1033:23:@1421.4]
  assign _T_2170 = _T_548[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:37:@1426.4]
  assign _T_2173 = _T_2002 <= 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:43:@1427.4]
  assign _T_2174 = _T_1998[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:87:@1428.4]
  assign _T_2176 = _T_2174 == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:91:@1429.4]
  assign _T_2177 = _T_2173 & _T_2176; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:72:@1430.4]
  assign _T_2179 = _T_2160[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:171:@1431.4]
  assign _T_2180 = {256'h0,_T_2179}; // @[Cat.scala 30:58:@1432.4]
  assign _T_2186 = _T_2173 & _T_2174; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:72:@1436.4]
  assign _T_2188 = _T_2160[511:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:171:@1437.4]
  assign _T_2189 = {256'h0,_T_2188}; // @[Cat.scala 30:58:@1438.4]
  assign _T_2190 = _T_2186 ? _T_2189 : _T_2160; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:27:@1439.4]
  assign _T_2191 = _T_2177 ? _T_2180 : _T_2190; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:27:@1440.4]
  assign _T_2192 = _T_2170 ? 512'h0 : _T_2191; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:27:@1441.4]
  assign _T_2263 = _T_2192[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1444.4]
  assign _T_2264 = _T_2192[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1446.4]
  assign _T_2265 = _T_2192[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1448.4]
  assign _T_2266 = _T_2192[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1450.4]
  assign _T_2267 = _T_2192[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1452.4]
  assign _T_2268 = _T_2192[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1454.4]
  assign _T_2269 = _T_2192[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1456.4]
  assign _T_2270 = _T_2192[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1458.4]
  assign _T_2271 = _T_2192[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1460.4]
  assign _T_2272 = _T_2192[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1462.4]
  assign _T_2273 = _T_2192[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1464.4]
  assign _T_2274 = _T_2192[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1466.4]
  assign _T_2275 = _T_2192[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1468.4]
  assign _T_2276 = _T_2192[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1470.4]
  assign _T_2277 = _T_2192[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1472.4]
  assign _T_2278 = _T_2192[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1474.4]
  assign _T_2279 = _T_2192[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1476.4]
  assign _T_2280 = _T_2192[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1478.4]
  assign _T_2281 = _T_2192[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1480.4]
  assign _T_2282 = _T_2192[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1482.4]
  assign _T_2283 = _T_2192[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1484.4]
  assign _T_2284 = _T_2192[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1486.4]
  assign _T_2285 = _T_2192[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1488.4]
  assign _T_2286 = _T_2192[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1490.4]
  assign _T_2287 = _T_2192[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1492.4]
  assign _T_2288 = _T_2192[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1494.4]
  assign _T_2289 = _T_2192[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1496.4]
  assign _T_2290 = _T_2192[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1498.4]
  assign _T_2291 = _T_2192[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1500.4]
  assign _T_2292 = _T_2192[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1502.4]
  assign _T_2293 = _T_2192[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1504.4]
  assign _T_2294 = _T_2192[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1506.4]
  assign _T_2295 = _T_2192[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1508.4]
  assign _T_2296 = _T_2192[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1510.4]
  assign _T_2297 = _T_2192[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1512.4]
  assign _T_2298 = _T_2192[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1514.4]
  assign _T_2299 = _T_2192[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1516.4]
  assign _T_2300 = _T_2192[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1518.4]
  assign _T_2301 = _T_2192[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1520.4]
  assign _T_2302 = _T_2192[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1522.4]
  assign _T_2303 = _T_2192[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1524.4]
  assign _T_2304 = _T_2192[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1526.4]
  assign _T_2305 = _T_2192[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1528.4]
  assign _T_2306 = _T_2192[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1530.4]
  assign _T_2307 = _T_2192[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1532.4]
  assign _T_2308 = _T_2192[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1534.4]
  assign _T_2309 = _T_2192[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1536.4]
  assign _T_2310 = _T_2192[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1538.4]
  assign _T_2311 = _T_2192[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1540.4]
  assign _T_2312 = _T_2192[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1542.4]
  assign _T_2313 = _T_2192[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1544.4]
  assign _T_2314 = _T_2192[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1546.4]
  assign _T_2315 = _T_2192[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1548.4]
  assign _T_2316 = _T_2192[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1550.4]
  assign _T_2317 = _T_2192[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1552.4]
  assign _T_2318 = _T_2192[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1554.4]
  assign _T_2319 = _T_2192[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1556.4]
  assign _T_2320 = _T_2192[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1558.4]
  assign _T_2321 = _T_2192[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1560.4]
  assign _T_2322 = _T_2192[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1562.4]
  assign _T_2323 = _T_2192[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1564.4]
  assign _T_2324 = _T_2192[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1566.4]
  assign _T_2325 = _T_2192[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1568.4]
  assign _T_2326 = _T_2192[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1570.4]
  assign _T_2339 = _T_548[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:39:@1578.4]
  assign _T_2340 = ~ _T_2339; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:29:@1579.4]
  assign _T_2342 = {_T_2160,_T_2164}; // @[Cat.scala 30:58:@1580.4]
  assign _T_2343 = _T_2340 ? 1024'h0 : _T_2342; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:28:@1581.4]
  assign _T_2344 = _T_548[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:39:@1582.4]
  assign _T_2345 = ~ _T_2344; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:29:@1583.4]
  assign _T_2347 = {_T_2158,_T_2158,_T_2158,_T_2158}; // @[Cat.scala 30:58:@1584.4]
  assign _T_2348 = _T_2345 ? 1024'h0 : _T_2347; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:28:@1585.4]
  assign _T_2349 = _T_548[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:39:@1586.4]
  assign _T_2350 = ~ _T_2349; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:29:@1587.4]
  assign _T_2353 = _T_2350 ? 1024'h0 : _T_2347; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:28:@1589.4]
  assign _T_2354 = _T_548[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:39:@1590.4]
  assign _T_2355 = ~ _T_2354; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:29:@1591.4]
  assign _T_2358 = _T_2355 ? 1024'h0 : _T_2347; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:28:@1593.4]
  assign _T_2360 = {_T_1899,3'h0}; // @[Cat.scala 30:58:@1594.4]
  assign _T_2361 = _T_2343 >> _T_2360; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:41:@1595.4]
  assign _T_2362 = _T_2361[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:82:@1596.4]
  assign _T_2364 = {_T_1902,3'h0}; // @[Cat.scala 30:58:@1597.4]
  assign _T_2365 = _T_2348 >> _T_2364; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:41:@1598.4]
  assign _T_2366 = _T_2365[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:82:@1599.4]
  assign _T_2368 = {_T_1905,3'h0}; // @[Cat.scala 30:58:@1600.4]
  assign _T_2369 = _T_2353 >> _T_2368; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:41:@1601.4]
  assign _T_2370 = _T_2369[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:82:@1602.4]
  assign _T_2372 = {_T_1908,3'h0}; // @[Cat.scala 30:58:@1603.4]
  assign _T_2373 = _T_2358 >> _T_2372; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:41:@1604.4]
  assign _T_2374 = _T_2373[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:82:@1605.4]
  assign _T_2375 = _T_548[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:36:@1606.4]
  assign _T_2376 = ~ _T_2375; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:26:@1607.4]
  assign _T_2379 = _T_610 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:41:@1608.4]
  assign _T_2380 = _T_2374[127:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:81:@1609.4]
  assign _T_2386 = {_T_2380,_T_2338,_T_2336,_T_2332}; // @[Cat.scala 30:58:@1615.4]
  assign _T_2388 = _T_610 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:41:@1616.4]
  assign _T_2389 = _T_2366[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:81:@1617.4]
  assign _T_2391 = {_T_2389,_T_2328}; // @[Cat.scala 30:58:@1619.4]
  assign _T_2393 = _T_2388 ? _T_2391 : _T_2362; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:25:@1621.4]
  assign _T_2394 = _T_2379 ? _T_2386 : _T_2393; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:25:@1622.4]
  assign _T_2395 = _T_2376 ? 512'h0 : _T_2394; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:25:@1623.4]
  assign _T_2466 = _T_2395[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1625.4]
  assign _T_2467 = _T_2395[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1627.4]
  assign _T_2468 = _T_2395[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1629.4]
  assign _T_2469 = _T_2395[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1631.4]
  assign _T_2470 = _T_2395[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1633.4]
  assign _T_2471 = _T_2395[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1635.4]
  assign _T_2472 = _T_2395[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1637.4]
  assign _T_2473 = _T_2395[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1639.4]
  assign _T_2474 = _T_2395[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1641.4]
  assign _T_2475 = _T_2395[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1643.4]
  assign _T_2476 = _T_2395[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1645.4]
  assign _T_2477 = _T_2395[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1647.4]
  assign _T_2478 = _T_2395[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1649.4]
  assign _T_2479 = _T_2395[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1651.4]
  assign _T_2480 = _T_2395[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1653.4]
  assign _T_2481 = _T_2395[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1655.4]
  assign _T_2482 = _T_2395[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1657.4]
  assign _T_2483 = _T_2395[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1659.4]
  assign _T_2484 = _T_2395[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1661.4]
  assign _T_2485 = _T_2395[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1663.4]
  assign _T_2486 = _T_2395[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1665.4]
  assign _T_2487 = _T_2395[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1667.4]
  assign _T_2488 = _T_2395[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1669.4]
  assign _T_2489 = _T_2395[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1671.4]
  assign _T_2490 = _T_2395[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1673.4]
  assign _T_2491 = _T_2395[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1675.4]
  assign _T_2492 = _T_2395[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1677.4]
  assign _T_2493 = _T_2395[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1679.4]
  assign _T_2494 = _T_2395[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1681.4]
  assign _T_2495 = _T_2395[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1683.4]
  assign _T_2496 = _T_2395[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1685.4]
  assign _T_2497 = _T_2395[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1687.4]
  assign _T_2498 = _T_2395[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1689.4]
  assign _T_2499 = _T_2395[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1691.4]
  assign _T_2500 = _T_2395[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1693.4]
  assign _T_2501 = _T_2395[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1695.4]
  assign _T_2502 = _T_2395[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1697.4]
  assign _T_2503 = _T_2395[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1699.4]
  assign _T_2504 = _T_2395[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1701.4]
  assign _T_2505 = _T_2395[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1703.4]
  assign _T_2506 = _T_2395[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1705.4]
  assign _T_2507 = _T_2395[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1707.4]
  assign _T_2508 = _T_2395[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1709.4]
  assign _T_2509 = _T_2395[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1711.4]
  assign _T_2510 = _T_2395[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1713.4]
  assign _T_2511 = _T_2395[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1715.4]
  assign _T_2512 = _T_2395[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1717.4]
  assign _T_2513 = _T_2395[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1719.4]
  assign _T_2514 = _T_2395[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1721.4]
  assign _T_2515 = _T_2395[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1723.4]
  assign _T_2516 = _T_2395[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1725.4]
  assign _T_2517 = _T_2395[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1727.4]
  assign _T_2518 = _T_2395[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1729.4]
  assign _T_2519 = _T_2395[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1731.4]
  assign _T_2520 = _T_2395[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1733.4]
  assign _T_2521 = _T_2395[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1735.4]
  assign _T_2522 = _T_2395[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1737.4]
  assign _T_2523 = _T_2395[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1739.4]
  assign _T_2524 = _T_2395[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1741.4]
  assign _T_2525 = _T_2395[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1743.4]
  assign _T_2526 = _T_2395[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1745.4]
  assign _T_2527 = _T_2395[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1747.4]
  assign _T_2528 = _T_2395[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1749.4]
  assign _T_2529 = _T_2395[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1751.4]
  assign _T_2531 = _T_613 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:59:@1753.4]
  assign _T_2532 = _T_1925 & _T_2531; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:41:@1754.4]
  assign _T_2534 = _T_613 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:59:@1755.4]
  assign _T_2535 = _T_1928 & _T_2534; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:41:@1756.4]
  assign _T_2538 = _T_1931 & _T_2534; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:41:@1758.4]
  assign _GEN_149 = _T_2532 ? _T_2362 : {{256'd0}, _T_2328}; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:24:@1759.4]
  assign _GEN_150 = _T_2535 ? _T_2328 : {{128'd0}, _T_2330}; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1762.4]
  assign _GEN_151 = _T_2535 ? _T_2366 : {{384'd0}, _T_2334}; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1762.4]
  assign _GEN_154 = _T_2538 ? _T_2370 : {{384'd0}, _T_2338}; // @[NV_NVDLA_CSC_dl_for_check.scala 1109:24:@1766.4]
  assign _T_2544 = 319'hffffffffffffffff << _T_2002; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:56:@1772.4]
  assign _T_2545 = _T_2544[63:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:73:@1773.4]
  assign _T_2546 = ~ _T_2545; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:24:@1774.4]
  assign _T_2548 = _T_2003 >= 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:51:@1775.4]
  assign _T_2555 = _T_2548 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:32:@1777.4]
  assign _T_2557 = _T_2003 >= 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:51:@1778.4]
  assign _T_2564 = _T_2557 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:32:@1780.4]
  assign _T_2566 = _T_2003 == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:51:@1781.4]
  assign _T_2573 = _T_2566 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:32:@1783.4]
  assign _T_2574 = _T_2555[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1124:57:@1784.4]
  assign _T_2580 = {_T_2574,32'hffffffff}; // @[Cat.scala 30:58:@1786.4]
  assign _T_2581 = _T_2573[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:57:@1787.4]
  assign _T_2582 = _T_2564[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:106:@1788.4]
  assign _T_2583 = _T_2555[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:155:@1789.4]
  assign _T_2591 = {_T_2581,_T_2582,_T_2583,16'hffff}; // @[Cat.scala 30:58:@1793.4]
  assign _T_2593 = _T_619 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:43:@1794.4]
  assign _T_2594 = _T_2546[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:89:@1795.4]
  assign _T_2596 = {_T_2594,_T_2594,_T_2594,_T_2594}; // @[Cat.scala 30:58:@1797.4]
  assign _T_2597 = _T_2596 & _T_2591; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:116:@1798.4]
  assign _T_2599 = _T_619 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:43:@1799.4]
  assign _T_2600 = _T_2546[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:89:@1800.4]
  assign _T_2601 = {_T_2600,_T_2600}; // @[Cat.scala 30:58:@1801.4]
  assign _T_2602 = _T_2601 & _T_2580; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:116:@1802.4]
  assign _T_2603 = _T_2599 ? _T_2602 : _T_2546; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:26:@1803.4]
  assign _T_2604 = _T_2593 ? _T_2597 : _T_2603; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:26:@1804.4]
  assign _T_2605 = _T_548[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:35:@1805.4]
  assign _T_2606_0 = _T_2605 ? _T_2466 : _T_2263; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_1 = _T_2605 ? _T_2467 : _T_2264; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_2 = _T_2605 ? _T_2468 : _T_2265; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_3 = _T_2605 ? _T_2469 : _T_2266; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_4 = _T_2605 ? _T_2470 : _T_2267; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_5 = _T_2605 ? _T_2471 : _T_2268; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_6 = _T_2605 ? _T_2472 : _T_2269; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_7 = _T_2605 ? _T_2473 : _T_2270; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_8 = _T_2605 ? _T_2474 : _T_2271; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_9 = _T_2605 ? _T_2475 : _T_2272; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_10 = _T_2605 ? _T_2476 : _T_2273; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_11 = _T_2605 ? _T_2477 : _T_2274; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_12 = _T_2605 ? _T_2478 : _T_2275; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_13 = _T_2605 ? _T_2479 : _T_2276; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_14 = _T_2605 ? _T_2480 : _T_2277; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_15 = _T_2605 ? _T_2481 : _T_2278; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_16 = _T_2605 ? _T_2482 : _T_2279; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_17 = _T_2605 ? _T_2483 : _T_2280; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_18 = _T_2605 ? _T_2484 : _T_2281; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_19 = _T_2605 ? _T_2485 : _T_2282; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_20 = _T_2605 ? _T_2486 : _T_2283; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_21 = _T_2605 ? _T_2487 : _T_2284; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_22 = _T_2605 ? _T_2488 : _T_2285; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_23 = _T_2605 ? _T_2489 : _T_2286; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_24 = _T_2605 ? _T_2490 : _T_2287; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_25 = _T_2605 ? _T_2491 : _T_2288; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_26 = _T_2605 ? _T_2492 : _T_2289; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_27 = _T_2605 ? _T_2493 : _T_2290; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_28 = _T_2605 ? _T_2494 : _T_2291; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_29 = _T_2605 ? _T_2495 : _T_2292; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_30 = _T_2605 ? _T_2496 : _T_2293; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_31 = _T_2605 ? _T_2497 : _T_2294; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_32 = _T_2605 ? _T_2498 : _T_2295; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_33 = _T_2605 ? _T_2499 : _T_2296; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_34 = _T_2605 ? _T_2500 : _T_2297; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_35 = _T_2605 ? _T_2501 : _T_2298; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_36 = _T_2605 ? _T_2502 : _T_2299; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_37 = _T_2605 ? _T_2503 : _T_2300; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_38 = _T_2605 ? _T_2504 : _T_2301; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_39 = _T_2605 ? _T_2505 : _T_2302; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_40 = _T_2605 ? _T_2506 : _T_2303; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_41 = _T_2605 ? _T_2507 : _T_2304; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_42 = _T_2605 ? _T_2508 : _T_2305; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_43 = _T_2605 ? _T_2509 : _T_2306; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_44 = _T_2605 ? _T_2510 : _T_2307; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_45 = _T_2605 ? _T_2511 : _T_2308; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_46 = _T_2605 ? _T_2512 : _T_2309; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_47 = _T_2605 ? _T_2513 : _T_2310; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_48 = _T_2605 ? _T_2514 : _T_2311; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_49 = _T_2605 ? _T_2515 : _T_2312; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_50 = _T_2605 ? _T_2516 : _T_2313; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_51 = _T_2605 ? _T_2517 : _T_2314; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_52 = _T_2605 ? _T_2518 : _T_2315; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_53 = _T_2605 ? _T_2519 : _T_2316; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_54 = _T_2605 ? _T_2520 : _T_2317; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_55 = _T_2605 ? _T_2521 : _T_2318; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_56 = _T_2605 ? _T_2522 : _T_2319; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_57 = _T_2605 ? _T_2523 : _T_2320; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_58 = _T_2605 ? _T_2524 : _T_2321; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_59 = _T_2605 ? _T_2525 : _T_2322; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_60 = _T_2605 ? _T_2526 : _T_2323; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_61 = _T_2605 ? _T_2527 : _T_2324; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_62 = _T_2605 ? _T_2528 : _T_2325; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2606_63 = _T_2605 ? _T_2529 : _T_2326; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1806.4]
  assign _T_2739 = _T_2606_0 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1807.4]
  assign _T_2741 = _T_2606_1 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1808.4]
  assign _T_2743 = _T_2606_2 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1809.4]
  assign _T_2745 = _T_2606_3 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1810.4]
  assign _T_2747 = _T_2606_4 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1811.4]
  assign _T_2749 = _T_2606_5 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1812.4]
  assign _T_2751 = _T_2606_6 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1813.4]
  assign _T_2753 = _T_2606_7 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1814.4]
  assign _T_2755 = _T_2606_8 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1815.4]
  assign _T_2757 = _T_2606_9 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1816.4]
  assign _T_2759 = _T_2606_10 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1817.4]
  assign _T_2761 = _T_2606_11 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1818.4]
  assign _T_2763 = _T_2606_12 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1819.4]
  assign _T_2765 = _T_2606_13 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1820.4]
  assign _T_2767 = _T_2606_14 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1821.4]
  assign _T_2769 = _T_2606_15 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1822.4]
  assign _T_2771 = _T_2606_16 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1823.4]
  assign _T_2773 = _T_2606_17 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1824.4]
  assign _T_2775 = _T_2606_18 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1825.4]
  assign _T_2777 = _T_2606_19 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1826.4]
  assign _T_2779 = _T_2606_20 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1827.4]
  assign _T_2781 = _T_2606_21 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1828.4]
  assign _T_2783 = _T_2606_22 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1829.4]
  assign _T_2785 = _T_2606_23 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1830.4]
  assign _T_2787 = _T_2606_24 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1831.4]
  assign _T_2789 = _T_2606_25 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1832.4]
  assign _T_2791 = _T_2606_26 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1833.4]
  assign _T_2793 = _T_2606_27 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1834.4]
  assign _T_2795 = _T_2606_28 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1835.4]
  assign _T_2797 = _T_2606_29 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1836.4]
  assign _T_2799 = _T_2606_30 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1837.4]
  assign _T_2801 = _T_2606_31 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1838.4]
  assign _T_2803 = _T_2606_32 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1839.4]
  assign _T_2805 = _T_2606_33 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1840.4]
  assign _T_2807 = _T_2606_34 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1841.4]
  assign _T_2809 = _T_2606_35 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1842.4]
  assign _T_2811 = _T_2606_36 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1843.4]
  assign _T_2813 = _T_2606_37 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1844.4]
  assign _T_2815 = _T_2606_38 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1845.4]
  assign _T_2817 = _T_2606_39 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1846.4]
  assign _T_2819 = _T_2606_40 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1847.4]
  assign _T_2821 = _T_2606_41 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1848.4]
  assign _T_2823 = _T_2606_42 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1849.4]
  assign _T_2825 = _T_2606_43 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1850.4]
  assign _T_2827 = _T_2606_44 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1851.4]
  assign _T_2829 = _T_2606_45 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1852.4]
  assign _T_2831 = _T_2606_46 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1853.4]
  assign _T_2833 = _T_2606_47 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1854.4]
  assign _T_2835 = _T_2606_48 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1855.4]
  assign _T_2837 = _T_2606_49 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1856.4]
  assign _T_2839 = _T_2606_50 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1857.4]
  assign _T_2841 = _T_2606_51 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1858.4]
  assign _T_2843 = _T_2606_52 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1859.4]
  assign _T_2845 = _T_2606_53 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1860.4]
  assign _T_2847 = _T_2606_54 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1861.4]
  assign _T_2849 = _T_2606_55 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1862.4]
  assign _T_2851 = _T_2606_56 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1863.4]
  assign _T_2853 = _T_2606_57 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1864.4]
  assign _T_2855 = _T_2606_58 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1865.4]
  assign _T_2857 = _T_2606_59 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1866.4]
  assign _T_2859 = _T_2606_60 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1867.4]
  assign _T_2861 = _T_2606_61 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1868.4]
  assign _T_2863 = _T_2606_62 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1869.4]
  assign _T_2865 = _T_2606_63 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1870.4]
  assign _T_2936 = _T_2604[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1936.4]
  assign _T_2937 = _T_2936 & _T_2739; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1937.4]
  assign _T_2938 = _T_2604[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1938.4]
  assign _T_2939 = _T_2938 & _T_2741; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1939.4]
  assign _T_2940 = _T_2604[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1940.4]
  assign _T_2941 = _T_2940 & _T_2743; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1941.4]
  assign _T_2942 = _T_2604[3]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1942.4]
  assign _T_2943 = _T_2942 & _T_2745; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1943.4]
  assign _T_2944 = _T_2604[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1944.4]
  assign _T_2945 = _T_2944 & _T_2747; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1945.4]
  assign _T_2946 = _T_2604[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1946.4]
  assign _T_2947 = _T_2946 & _T_2749; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1947.4]
  assign _T_2948 = _T_2604[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1948.4]
  assign _T_2949 = _T_2948 & _T_2751; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1949.4]
  assign _T_2950 = _T_2604[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1950.4]
  assign _T_2951 = _T_2950 & _T_2753; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1951.4]
  assign _T_2952 = _T_2604[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1952.4]
  assign _T_2953 = _T_2952 & _T_2755; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1953.4]
  assign _T_2954 = _T_2604[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1954.4]
  assign _T_2955 = _T_2954 & _T_2757; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1955.4]
  assign _T_2956 = _T_2604[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1956.4]
  assign _T_2957 = _T_2956 & _T_2759; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1957.4]
  assign _T_2958 = _T_2604[11]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1958.4]
  assign _T_2959 = _T_2958 & _T_2761; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1959.4]
  assign _T_2960 = _T_2604[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1960.4]
  assign _T_2961 = _T_2960 & _T_2763; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1961.4]
  assign _T_2962 = _T_2604[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1962.4]
  assign _T_2963 = _T_2962 & _T_2765; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1963.4]
  assign _T_2964 = _T_2604[14]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1964.4]
  assign _T_2965 = _T_2964 & _T_2767; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1965.4]
  assign _T_2966 = _T_2604[15]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1966.4]
  assign _T_2967 = _T_2966 & _T_2769; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1967.4]
  assign _T_2968 = _T_2604[16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1968.4]
  assign _T_2969 = _T_2968 & _T_2771; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1969.4]
  assign _T_2970 = _T_2604[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1970.4]
  assign _T_2971 = _T_2970 & _T_2773; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1971.4]
  assign _T_2972 = _T_2604[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1972.4]
  assign _T_2973 = _T_2972 & _T_2775; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1973.4]
  assign _T_2974 = _T_2604[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1974.4]
  assign _T_2975 = _T_2974 & _T_2777; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1975.4]
  assign _T_2976 = _T_2604[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1976.4]
  assign _T_2977 = _T_2976 & _T_2779; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1977.4]
  assign _T_2978 = _T_2604[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1978.4]
  assign _T_2979 = _T_2978 & _T_2781; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1979.4]
  assign _T_2980 = _T_2604[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1980.4]
  assign _T_2981 = _T_2980 & _T_2783; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1981.4]
  assign _T_2982 = _T_2604[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1982.4]
  assign _T_2983 = _T_2982 & _T_2785; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1983.4]
  assign _T_2984 = _T_2604[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1984.4]
  assign _T_2985 = _T_2984 & _T_2787; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1985.4]
  assign _T_2986 = _T_2604[25]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1986.4]
  assign _T_2987 = _T_2986 & _T_2789; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1987.4]
  assign _T_2988 = _T_2604[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1988.4]
  assign _T_2989 = _T_2988 & _T_2791; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1989.4]
  assign _T_2990 = _T_2604[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1990.4]
  assign _T_2991 = _T_2990 & _T_2793; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1991.4]
  assign _T_2992 = _T_2604[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1992.4]
  assign _T_2993 = _T_2992 & _T_2795; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1993.4]
  assign _T_2994 = _T_2604[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1994.4]
  assign _T_2995 = _T_2994 & _T_2797; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1995.4]
  assign _T_2996 = _T_2604[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1996.4]
  assign _T_2997 = _T_2996 & _T_2799; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1997.4]
  assign _T_2998 = _T_2604[31]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1998.4]
  assign _T_2999 = _T_2998 & _T_2801; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1999.4]
  assign _T_3000 = _T_2604[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2000.4]
  assign _T_3001 = _T_3000 & _T_2803; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2001.4]
  assign _T_3002 = _T_2604[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2002.4]
  assign _T_3003 = _T_3002 & _T_2805; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2003.4]
  assign _T_3004 = _T_2604[34]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2004.4]
  assign _T_3005 = _T_3004 & _T_2807; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2005.4]
  assign _T_3006 = _T_2604[35]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2006.4]
  assign _T_3007 = _T_3006 & _T_2809; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2007.4]
  assign _T_3008 = _T_2604[36]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2008.4]
  assign _T_3009 = _T_3008 & _T_2811; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2009.4]
  assign _T_3010 = _T_2604[37]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2010.4]
  assign _T_3011 = _T_3010 & _T_2813; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2011.4]
  assign _T_3012 = _T_2604[38]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2012.4]
  assign _T_3013 = _T_3012 & _T_2815; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2013.4]
  assign _T_3014 = _T_2604[39]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2014.4]
  assign _T_3015 = _T_3014 & _T_2817; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2015.4]
  assign _T_3016 = _T_2604[40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2016.4]
  assign _T_3017 = _T_3016 & _T_2819; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2017.4]
  assign _T_3018 = _T_2604[41]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2018.4]
  assign _T_3019 = _T_3018 & _T_2821; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2019.4]
  assign _T_3020 = _T_2604[42]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2020.4]
  assign _T_3021 = _T_3020 & _T_2823; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2021.4]
  assign _T_3022 = _T_2604[43]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2022.4]
  assign _T_3023 = _T_3022 & _T_2825; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2023.4]
  assign _T_3024 = _T_2604[44]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2024.4]
  assign _T_3025 = _T_3024 & _T_2827; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2025.4]
  assign _T_3026 = _T_2604[45]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2026.4]
  assign _T_3027 = _T_3026 & _T_2829; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2027.4]
  assign _T_3028 = _T_2604[46]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2028.4]
  assign _T_3029 = _T_3028 & _T_2831; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2029.4]
  assign _T_3030 = _T_2604[47]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2030.4]
  assign _T_3031 = _T_3030 & _T_2833; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2031.4]
  assign _T_3032 = _T_2604[48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2032.4]
  assign _T_3033 = _T_3032 & _T_2835; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2033.4]
  assign _T_3034 = _T_2604[49]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2034.4]
  assign _T_3035 = _T_3034 & _T_2837; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2035.4]
  assign _T_3036 = _T_2604[50]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2036.4]
  assign _T_3037 = _T_3036 & _T_2839; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2037.4]
  assign _T_3038 = _T_2604[51]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2038.4]
  assign _T_3039 = _T_3038 & _T_2841; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2039.4]
  assign _T_3040 = _T_2604[52]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2040.4]
  assign _T_3041 = _T_3040 & _T_2843; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2041.4]
  assign _T_3042 = _T_2604[53]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2042.4]
  assign _T_3043 = _T_3042 & _T_2845; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2043.4]
  assign _T_3044 = _T_2604[54]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2044.4]
  assign _T_3045 = _T_3044 & _T_2847; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2045.4]
  assign _T_3046 = _T_2604[55]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2046.4]
  assign _T_3047 = _T_3046 & _T_2849; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2047.4]
  assign _T_3048 = _T_2604[56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2048.4]
  assign _T_3049 = _T_3048 & _T_2851; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2049.4]
  assign _T_3050 = _T_2604[57]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2050.4]
  assign _T_3051 = _T_3050 & _T_2853; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2051.4]
  assign _T_3052 = _T_2604[58]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2052.4]
  assign _T_3053 = _T_3052 & _T_2855; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2053.4]
  assign _T_3054 = _T_2604[59]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2054.4]
  assign _T_3055 = _T_3054 & _T_2857; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2055.4]
  assign _T_3056 = _T_2604[60]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2056.4]
  assign _T_3057 = _T_3056 & _T_2859; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2057.4]
  assign _T_3058 = _T_2604[61]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2058.4]
  assign _T_3059 = _T_3058 & _T_2861; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2059.4]
  assign _T_3060 = _T_2604[62]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2060.4]
  assign _T_3061 = _T_3060 & _T_2863; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2061.4]
  assign _T_3062 = _T_2604[63]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2062.4]
  assign _T_3063 = _T_3062 & _T_2865; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2063.4]
  assign _GEN_156 = _T_1965 ? _T_2937 : _T_3406_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_157 = _T_1965 ? _T_2939 : _T_3406_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_158 = _T_1965 ? _T_2941 : _T_3406_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_159 = _T_1965 ? _T_2943 : _T_3406_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_160 = _T_1965 ? _T_2945 : _T_3406_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_161 = _T_1965 ? _T_2947 : _T_3406_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_162 = _T_1965 ? _T_2949 : _T_3406_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_163 = _T_1965 ? _T_2951 : _T_3406_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_164 = _T_1965 ? _T_2953 : _T_3406_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_165 = _T_1965 ? _T_2955 : _T_3406_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_166 = _T_1965 ? _T_2957 : _T_3406_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_167 = _T_1965 ? _T_2959 : _T_3406_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_168 = _T_1965 ? _T_2961 : _T_3406_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_169 = _T_1965 ? _T_2963 : _T_3406_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_170 = _T_1965 ? _T_2965 : _T_3406_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_171 = _T_1965 ? _T_2967 : _T_3406_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_172 = _T_1965 ? _T_2969 : _T_3406_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_173 = _T_1965 ? _T_2971 : _T_3406_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_174 = _T_1965 ? _T_2973 : _T_3406_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_175 = _T_1965 ? _T_2975 : _T_3406_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_176 = _T_1965 ? _T_2977 : _T_3406_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_177 = _T_1965 ? _T_2979 : _T_3406_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_178 = _T_1965 ? _T_2981 : _T_3406_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_179 = _T_1965 ? _T_2983 : _T_3406_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_180 = _T_1965 ? _T_2985 : _T_3406_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_181 = _T_1965 ? _T_2987 : _T_3406_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_182 = _T_1965 ? _T_2989 : _T_3406_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_183 = _T_1965 ? _T_2991 : _T_3406_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_184 = _T_1965 ? _T_2993 : _T_3406_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_185 = _T_1965 ? _T_2995 : _T_3406_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_186 = _T_1965 ? _T_2997 : _T_3406_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_187 = _T_1965 ? _T_2999 : _T_3406_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_188 = _T_1965 ? _T_3001 : _T_3406_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_189 = _T_1965 ? _T_3003 : _T_3406_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_190 = _T_1965 ? _T_3005 : _T_3406_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_191 = _T_1965 ? _T_3007 : _T_3406_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_192 = _T_1965 ? _T_3009 : _T_3406_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_193 = _T_1965 ? _T_3011 : _T_3406_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_194 = _T_1965 ? _T_3013 : _T_3406_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_195 = _T_1965 ? _T_3015 : _T_3406_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_196 = _T_1965 ? _T_3017 : _T_3406_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_197 = _T_1965 ? _T_3019 : _T_3406_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_198 = _T_1965 ? _T_3021 : _T_3406_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_199 = _T_1965 ? _T_3023 : _T_3406_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_200 = _T_1965 ? _T_3025 : _T_3406_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_201 = _T_1965 ? _T_3027 : _T_3406_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_202 = _T_1965 ? _T_3029 : _T_3406_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_203 = _T_1965 ? _T_3031 : _T_3406_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_204 = _T_1965 ? _T_3033 : _T_3406_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_205 = _T_1965 ? _T_3035 : _T_3406_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_206 = _T_1965 ? _T_3037 : _T_3406_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_207 = _T_1965 ? _T_3039 : _T_3406_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_208 = _T_1965 ? _T_3041 : _T_3406_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_209 = _T_1965 ? _T_3043 : _T_3406_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_210 = _T_1965 ? _T_3045 : _T_3406_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_211 = _T_1965 ? _T_3047 : _T_3406_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_212 = _T_1965 ? _T_3049 : _T_3406_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_213 = _T_1965 ? _T_3051 : _T_3406_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_214 = _T_1965 ? _T_3053 : _T_3406_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_215 = _T_1965 ? _T_3055 : _T_3406_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_216 = _T_1965 ? _T_3057 : _T_3406_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_217 = _T_1965 ? _T_3059 : _T_3406_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_218 = _T_1965 ? _T_3061 : _T_3406_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _GEN_219 = _T_1965 ? _T_3063 : _T_3406_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2202.4]
  assign _T_3673 = _T_1965 & _T_2937; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2268.4]
  assign _T_3674 = _T_1965 & _T_2939; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2272.4]
  assign _T_3675 = _T_1965 & _T_2941; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2276.4]
  assign _T_3676 = _T_1965 & _T_2943; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2280.4]
  assign _T_3677 = _T_1965 & _T_2945; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2284.4]
  assign _T_3678 = _T_1965 & _T_2947; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2288.4]
  assign _T_3679 = _T_1965 & _T_2949; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2292.4]
  assign _T_3680 = _T_1965 & _T_2951; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2296.4]
  assign _T_3681 = _T_1965 & _T_2953; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2300.4]
  assign _T_3682 = _T_1965 & _T_2955; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2304.4]
  assign _T_3683 = _T_1965 & _T_2957; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2308.4]
  assign _T_3684 = _T_1965 & _T_2959; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2312.4]
  assign _T_3685 = _T_1965 & _T_2961; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2316.4]
  assign _T_3686 = _T_1965 & _T_2963; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2320.4]
  assign _T_3687 = _T_1965 & _T_2965; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2324.4]
  assign _T_3688 = _T_1965 & _T_2967; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2328.4]
  assign _T_3689 = _T_1965 & _T_2969; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2332.4]
  assign _T_3690 = _T_1965 & _T_2971; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2336.4]
  assign _T_3691 = _T_1965 & _T_2973; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2340.4]
  assign _T_3692 = _T_1965 & _T_2975; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2344.4]
  assign _T_3693 = _T_1965 & _T_2977; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2348.4]
  assign _T_3694 = _T_1965 & _T_2979; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2352.4]
  assign _T_3695 = _T_1965 & _T_2981; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2356.4]
  assign _T_3696 = _T_1965 & _T_2983; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2360.4]
  assign _T_3697 = _T_1965 & _T_2985; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2364.4]
  assign _T_3698 = _T_1965 & _T_2987; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2368.4]
  assign _T_3699 = _T_1965 & _T_2989; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2372.4]
  assign _T_3700 = _T_1965 & _T_2991; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2376.4]
  assign _T_3701 = _T_1965 & _T_2993; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2380.4]
  assign _T_3702 = _T_1965 & _T_2995; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2384.4]
  assign _T_3703 = _T_1965 & _T_2997; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2388.4]
  assign _T_3704 = _T_1965 & _T_2999; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2392.4]
  assign _T_3705 = _T_1965 & _T_3001; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2396.4]
  assign _T_3706 = _T_1965 & _T_3003; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2400.4]
  assign _T_3707 = _T_1965 & _T_3005; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2404.4]
  assign _T_3708 = _T_1965 & _T_3007; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2408.4]
  assign _T_3709 = _T_1965 & _T_3009; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2412.4]
  assign _T_3710 = _T_1965 & _T_3011; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2416.4]
  assign _T_3711 = _T_1965 & _T_3013; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2420.4]
  assign _T_3712 = _T_1965 & _T_3015; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2424.4]
  assign _T_3713 = _T_1965 & _T_3017; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2428.4]
  assign _T_3714 = _T_1965 & _T_3019; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2432.4]
  assign _T_3715 = _T_1965 & _T_3021; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2436.4]
  assign _T_3716 = _T_1965 & _T_3023; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2440.4]
  assign _T_3717 = _T_1965 & _T_3025; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2444.4]
  assign _T_3718 = _T_1965 & _T_3027; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2448.4]
  assign _T_3719 = _T_1965 & _T_3029; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2452.4]
  assign _T_3720 = _T_1965 & _T_3031; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2456.4]
  assign _T_3721 = _T_1965 & _T_3033; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2460.4]
  assign _T_3722 = _T_1965 & _T_3035; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2464.4]
  assign _T_3723 = _T_1965 & _T_3037; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2468.4]
  assign _T_3724 = _T_1965 & _T_3039; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2472.4]
  assign _T_3725 = _T_1965 & _T_3041; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2476.4]
  assign _T_3726 = _T_1965 & _T_3043; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2480.4]
  assign _T_3727 = _T_1965 & _T_3045; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2484.4]
  assign _T_3728 = _T_1965 & _T_3047; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2488.4]
  assign _T_3729 = _T_1965 & _T_3049; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2492.4]
  assign _T_3730 = _T_1965 & _T_3051; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2496.4]
  assign _T_3731 = _T_1965 & _T_3053; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2500.4]
  assign _T_3732 = _T_1965 & _T_3055; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2504.4]
  assign _T_3733 = _T_1965 & _T_3057; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2508.4]
  assign _T_3734 = _T_1965 & _T_3059; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2512.4]
  assign _T_3735 = _T_1965 & _T_3061; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2516.4]
  assign _T_3736 = _T_1965 & _T_3063; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2520.4]
  assign _T_4276 = ~ _T_3136; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:24:@2593.4]
  assign _T_4411_0 = _T_4276 ? 1'h0 : _T_3406_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_1 = _T_4276 ? 1'h0 : _T_3406_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_2 = _T_4276 ? 1'h0 : _T_3406_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_3 = _T_4276 ? 1'h0 : _T_3406_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_4 = _T_4276 ? 1'h0 : _T_3406_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_5 = _T_4276 ? 1'h0 : _T_3406_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_6 = _T_4276 ? 1'h0 : _T_3406_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_7 = _T_4276 ? 1'h0 : _T_3406_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_8 = _T_4276 ? 1'h0 : _T_3406_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_9 = _T_4276 ? 1'h0 : _T_3406_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_10 = _T_4276 ? 1'h0 : _T_3406_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_11 = _T_4276 ? 1'h0 : _T_3406_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_12 = _T_4276 ? 1'h0 : _T_3406_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_13 = _T_4276 ? 1'h0 : _T_3406_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_14 = _T_4276 ? 1'h0 : _T_3406_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_15 = _T_4276 ? 1'h0 : _T_3406_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_16 = _T_4276 ? 1'h0 : _T_3406_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_17 = _T_4276 ? 1'h0 : _T_3406_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_18 = _T_4276 ? 1'h0 : _T_3406_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_19 = _T_4276 ? 1'h0 : _T_3406_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_20 = _T_4276 ? 1'h0 : _T_3406_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_21 = _T_4276 ? 1'h0 : _T_3406_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_22 = _T_4276 ? 1'h0 : _T_3406_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_23 = _T_4276 ? 1'h0 : _T_3406_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_24 = _T_4276 ? 1'h0 : _T_3406_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_25 = _T_4276 ? 1'h0 : _T_3406_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_26 = _T_4276 ? 1'h0 : _T_3406_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_27 = _T_4276 ? 1'h0 : _T_3406_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_28 = _T_4276 ? 1'h0 : _T_3406_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_29 = _T_4276 ? 1'h0 : _T_3406_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_30 = _T_4276 ? 1'h0 : _T_3406_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_31 = _T_4276 ? 1'h0 : _T_3406_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_32 = _T_4276 ? 1'h0 : _T_3406_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_33 = _T_4276 ? 1'h0 : _T_3406_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_34 = _T_4276 ? 1'h0 : _T_3406_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_35 = _T_4276 ? 1'h0 : _T_3406_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_36 = _T_4276 ? 1'h0 : _T_3406_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_37 = _T_4276 ? 1'h0 : _T_3406_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_38 = _T_4276 ? 1'h0 : _T_3406_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_39 = _T_4276 ? 1'h0 : _T_3406_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_40 = _T_4276 ? 1'h0 : _T_3406_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_41 = _T_4276 ? 1'h0 : _T_3406_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_42 = _T_4276 ? 1'h0 : _T_3406_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_43 = _T_4276 ? 1'h0 : _T_3406_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_44 = _T_4276 ? 1'h0 : _T_3406_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_45 = _T_4276 ? 1'h0 : _T_3406_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_46 = _T_4276 ? 1'h0 : _T_3406_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_47 = _T_4276 ? 1'h0 : _T_3406_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_48 = _T_4276 ? 1'h0 : _T_3406_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_49 = _T_4276 ? 1'h0 : _T_3406_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_50 = _T_4276 ? 1'h0 : _T_3406_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_51 = _T_4276 ? 1'h0 : _T_3406_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_52 = _T_4276 ? 1'h0 : _T_3406_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_53 = _T_4276 ? 1'h0 : _T_3406_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_54 = _T_4276 ? 1'h0 : _T_3406_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_55 = _T_4276 ? 1'h0 : _T_3406_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_56 = _T_4276 ? 1'h0 : _T_3406_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_57 = _T_4276 ? 1'h0 : _T_3406_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_58 = _T_4276 ? 1'h0 : _T_3406_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_59 = _T_4276 ? 1'h0 : _T_3406_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_60 = _T_4276 ? 1'h0 : _T_3406_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_61 = _T_4276 ? 1'h0 : _T_3406_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_62 = _T_4276 ? 1'h0 : _T_3406_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4411_63 = _T_4276 ? 1'h0 : _T_3406_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2659.4]
  assign _T_4543 = _T_3136 | _T_3739; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:19:@2661.4]
  assign _GEN_284 = _T_4543 ? _T_4411_0 : _T_4006_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_285 = _T_4543 ? _T_4411_1 : _T_4006_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_286 = _T_4543 ? _T_4411_2 : _T_4006_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_287 = _T_4543 ? _T_4411_3 : _T_4006_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_288 = _T_4543 ? _T_4411_4 : _T_4006_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_289 = _T_4543 ? _T_4411_5 : _T_4006_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_290 = _T_4543 ? _T_4411_6 : _T_4006_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_291 = _T_4543 ? _T_4411_7 : _T_4006_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_292 = _T_4543 ? _T_4411_8 : _T_4006_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_293 = _T_4543 ? _T_4411_9 : _T_4006_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_294 = _T_4543 ? _T_4411_10 : _T_4006_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_295 = _T_4543 ? _T_4411_11 : _T_4006_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_296 = _T_4543 ? _T_4411_12 : _T_4006_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_297 = _T_4543 ? _T_4411_13 : _T_4006_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_298 = _T_4543 ? _T_4411_14 : _T_4006_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_299 = _T_4543 ? _T_4411_15 : _T_4006_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_300 = _T_4543 ? _T_4411_16 : _T_4006_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_301 = _T_4543 ? _T_4411_17 : _T_4006_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_302 = _T_4543 ? _T_4411_18 : _T_4006_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_303 = _T_4543 ? _T_4411_19 : _T_4006_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_304 = _T_4543 ? _T_4411_20 : _T_4006_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_305 = _T_4543 ? _T_4411_21 : _T_4006_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_306 = _T_4543 ? _T_4411_22 : _T_4006_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_307 = _T_4543 ? _T_4411_23 : _T_4006_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_308 = _T_4543 ? _T_4411_24 : _T_4006_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_309 = _T_4543 ? _T_4411_25 : _T_4006_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_310 = _T_4543 ? _T_4411_26 : _T_4006_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_311 = _T_4543 ? _T_4411_27 : _T_4006_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_312 = _T_4543 ? _T_4411_28 : _T_4006_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_313 = _T_4543 ? _T_4411_29 : _T_4006_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_314 = _T_4543 ? _T_4411_30 : _T_4006_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_315 = _T_4543 ? _T_4411_31 : _T_4006_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_316 = _T_4543 ? _T_4411_32 : _T_4006_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_317 = _T_4543 ? _T_4411_33 : _T_4006_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_318 = _T_4543 ? _T_4411_34 : _T_4006_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_319 = _T_4543 ? _T_4411_35 : _T_4006_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_320 = _T_4543 ? _T_4411_36 : _T_4006_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_321 = _T_4543 ? _T_4411_37 : _T_4006_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_322 = _T_4543 ? _T_4411_38 : _T_4006_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_323 = _T_4543 ? _T_4411_39 : _T_4006_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_324 = _T_4543 ? _T_4411_40 : _T_4006_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_325 = _T_4543 ? _T_4411_41 : _T_4006_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_326 = _T_4543 ? _T_4411_42 : _T_4006_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_327 = _T_4543 ? _T_4411_43 : _T_4006_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_328 = _T_4543 ? _T_4411_44 : _T_4006_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_329 = _T_4543 ? _T_4411_45 : _T_4006_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_330 = _T_4543 ? _T_4411_46 : _T_4006_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_331 = _T_4543 ? _T_4411_47 : _T_4006_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_332 = _T_4543 ? _T_4411_48 : _T_4006_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_333 = _T_4543 ? _T_4411_49 : _T_4006_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_334 = _T_4543 ? _T_4411_50 : _T_4006_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_335 = _T_4543 ? _T_4411_51 : _T_4006_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_336 = _T_4543 ? _T_4411_52 : _T_4006_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_337 = _T_4543 ? _T_4411_53 : _T_4006_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_338 = _T_4543 ? _T_4411_54 : _T_4006_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_339 = _T_4543 ? _T_4411_55 : _T_4006_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_340 = _T_4543 ? _T_4411_56 : _T_4006_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_341 = _T_4543 ? _T_4411_57 : _T_4006_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_342 = _T_4543 ? _T_4411_58 : _T_4006_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_343 = _T_4543 ? _T_4411_59 : _T_4006_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_344 = _T_4543 ? _T_4411_60 : _T_4006_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_345 = _T_4543 ? _T_4411_61 : _T_4006_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_346 = _T_4543 ? _T_4411_62 : _T_4006_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_347 = _T_4543 ? _T_4411_63 : _T_4006_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2662.4]
  assign _GEN_348 = _T_3136 ? {{8'd0}, _T_3136} : _T_4205; // @[NV_NVDLA_CSC_dl_for_check.scala 1182:19:@2728.4]
  assign _T_4547 = ~ _T_3739; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:27:@2925.4]
  assign _T_4549 = _T_4547 ? 9'h0 : _T_4205; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:26:@2926.4]
  assign _T_4557 = _T_3739 | _T_4546; // @[NV_NVDLA_CSC_dl_for_check.scala 1200:85:@2933.4]
  assign _GEN_413 = _T_4557 ? _T_4549 : _T_4559; // @[Reg.scala 20:19:@2935.4]
  assign _GEN_414 = _T_4557 ? _T_4549 : _T_4563; // @[Reg.scala 20:19:@2941.4]
  assign _GEN_415 = _T_4557 ? _T_4006_0 : _T_4831_0; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_416 = _T_4557 ? _T_4006_1 : _T_4831_1; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_417 = _T_4557 ? _T_4006_2 : _T_4831_2; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_418 = _T_4557 ? _T_4006_3 : _T_4831_3; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_419 = _T_4557 ? _T_4006_4 : _T_4831_4; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_420 = _T_4557 ? _T_4006_5 : _T_4831_5; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_421 = _T_4557 ? _T_4006_6 : _T_4831_6; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_422 = _T_4557 ? _T_4006_7 : _T_4831_7; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_423 = _T_4557 ? _T_4006_8 : _T_4831_8; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_424 = _T_4557 ? _T_4006_9 : _T_4831_9; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_425 = _T_4557 ? _T_4006_10 : _T_4831_10; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_426 = _T_4557 ? _T_4006_11 : _T_4831_11; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_427 = _T_4557 ? _T_4006_12 : _T_4831_12; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_428 = _T_4557 ? _T_4006_13 : _T_4831_13; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_429 = _T_4557 ? _T_4006_14 : _T_4831_14; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_430 = _T_4557 ? _T_4006_15 : _T_4831_15; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_431 = _T_4557 ? _T_4006_16 : _T_4831_16; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_432 = _T_4557 ? _T_4006_17 : _T_4831_17; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_433 = _T_4557 ? _T_4006_18 : _T_4831_18; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_434 = _T_4557 ? _T_4006_19 : _T_4831_19; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_435 = _T_4557 ? _T_4006_20 : _T_4831_20; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_436 = _T_4557 ? _T_4006_21 : _T_4831_21; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_437 = _T_4557 ? _T_4006_22 : _T_4831_22; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_438 = _T_4557 ? _T_4006_23 : _T_4831_23; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_439 = _T_4557 ? _T_4006_24 : _T_4831_24; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_440 = _T_4557 ? _T_4006_25 : _T_4831_25; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_441 = _T_4557 ? _T_4006_26 : _T_4831_26; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_442 = _T_4557 ? _T_4006_27 : _T_4831_27; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_443 = _T_4557 ? _T_4006_28 : _T_4831_28; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_444 = _T_4557 ? _T_4006_29 : _T_4831_29; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_445 = _T_4557 ? _T_4006_30 : _T_4831_30; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_446 = _T_4557 ? _T_4006_31 : _T_4831_31; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_447 = _T_4557 ? _T_4006_32 : _T_4831_32; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_448 = _T_4557 ? _T_4006_33 : _T_4831_33; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_449 = _T_4557 ? _T_4006_34 : _T_4831_34; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_450 = _T_4557 ? _T_4006_35 : _T_4831_35; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_451 = _T_4557 ? _T_4006_36 : _T_4831_36; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_452 = _T_4557 ? _T_4006_37 : _T_4831_37; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_453 = _T_4557 ? _T_4006_38 : _T_4831_38; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_454 = _T_4557 ? _T_4006_39 : _T_4831_39; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_455 = _T_4557 ? _T_4006_40 : _T_4831_40; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_456 = _T_4557 ? _T_4006_41 : _T_4831_41; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_457 = _T_4557 ? _T_4006_42 : _T_4831_42; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_458 = _T_4557 ? _T_4006_43 : _T_4831_43; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_459 = _T_4557 ? _T_4006_44 : _T_4831_44; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_460 = _T_4557 ? _T_4006_45 : _T_4831_45; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_461 = _T_4557 ? _T_4006_46 : _T_4831_46; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_462 = _T_4557 ? _T_4006_47 : _T_4831_47; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_463 = _T_4557 ? _T_4006_48 : _T_4831_48; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_464 = _T_4557 ? _T_4006_49 : _T_4831_49; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_465 = _T_4557 ? _T_4006_50 : _T_4831_50; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_466 = _T_4557 ? _T_4006_51 : _T_4831_51; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_467 = _T_4557 ? _T_4006_52 : _T_4831_52; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_468 = _T_4557 ? _T_4006_53 : _T_4831_53; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_469 = _T_4557 ? _T_4006_54 : _T_4831_54; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_470 = _T_4557 ? _T_4006_55 : _T_4831_55; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_471 = _T_4557 ? _T_4006_56 : _T_4831_56; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_472 = _T_4557 ? _T_4006_57 : _T_4831_57; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_473 = _T_4557 ? _T_4006_58 : _T_4831_58; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_474 = _T_4557 ? _T_4006_59 : _T_4831_59; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_475 = _T_4557 ? _T_4006_60 : _T_4831_60; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_476 = _T_4557 ? _T_4006_61 : _T_4831_61; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_477 = _T_4557 ? _T_4006_62 : _T_4831_62; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_478 = _T_4557 ? _T_4006_63 : _T_4831_63; // @[Reg.scala 20:19:@3012.4]
  assign _T_5034 = {_T_4831_7,_T_4831_6,_T_4831_5,_T_4831_4,_T_4831_3,_T_4831_2,_T_4831_1,_T_4831_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3084.4]
  assign _T_5042 = {_T_4831_15,_T_4831_14,_T_4831_13,_T_4831_12,_T_4831_11,_T_4831_10,_T_4831_9,_T_4831_8,_T_5034}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3092.4]
  assign _T_5049 = {_T_4831_23,_T_4831_22,_T_4831_21,_T_4831_20,_T_4831_19,_T_4831_18,_T_4831_17,_T_4831_16}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3099.4]
  assign _T_5058 = {_T_4831_31,_T_4831_30,_T_4831_29,_T_4831_28,_T_4831_27,_T_4831_26,_T_4831_25,_T_4831_24,_T_5049,_T_5042}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3108.4]
  assign _T_5065 = {_T_4831_39,_T_4831_38,_T_4831_37,_T_4831_36,_T_4831_35,_T_4831_34,_T_4831_33,_T_4831_32}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3115.4]
  assign _T_5073 = {_T_4831_47,_T_4831_46,_T_4831_45,_T_4831_44,_T_4831_43,_T_4831_42,_T_4831_41,_T_4831_40,_T_5065}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3123.4]
  assign _T_5080 = {_T_4831_55,_T_4831_54,_T_4831_53,_T_4831_52,_T_4831_51,_T_4831_50,_T_4831_49,_T_4831_48}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3130.4]
  assign _T_5089 = {_T_4831_63,_T_4831_62,_T_4831_61,_T_4831_60,_T_4831_59,_T_4831_58,_T_4831_57,_T_4831_56,_T_5080,_T_5073}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3139.4]
  assign _GEN_479 = _T_4557 ? _T_4006_0 : _T_5358_0; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_480 = _T_4557 ? _T_4006_1 : _T_5358_1; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_481 = _T_4557 ? _T_4006_2 : _T_5358_2; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_482 = _T_4557 ? _T_4006_3 : _T_5358_3; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_483 = _T_4557 ? _T_4006_4 : _T_5358_4; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_484 = _T_4557 ? _T_4006_5 : _T_5358_5; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_485 = _T_4557 ? _T_4006_6 : _T_5358_6; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_486 = _T_4557 ? _T_4006_7 : _T_5358_7; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_487 = _T_4557 ? _T_4006_8 : _T_5358_8; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_488 = _T_4557 ? _T_4006_9 : _T_5358_9; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_489 = _T_4557 ? _T_4006_10 : _T_5358_10; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_490 = _T_4557 ? _T_4006_11 : _T_5358_11; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_491 = _T_4557 ? _T_4006_12 : _T_5358_12; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_492 = _T_4557 ? _T_4006_13 : _T_5358_13; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_493 = _T_4557 ? _T_4006_14 : _T_5358_14; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_494 = _T_4557 ? _T_4006_15 : _T_5358_15; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_495 = _T_4557 ? _T_4006_16 : _T_5358_16; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_496 = _T_4557 ? _T_4006_17 : _T_5358_17; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_497 = _T_4557 ? _T_4006_18 : _T_5358_18; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_498 = _T_4557 ? _T_4006_19 : _T_5358_19; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_499 = _T_4557 ? _T_4006_20 : _T_5358_20; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_500 = _T_4557 ? _T_4006_21 : _T_5358_21; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_501 = _T_4557 ? _T_4006_22 : _T_5358_22; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_502 = _T_4557 ? _T_4006_23 : _T_5358_23; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_503 = _T_4557 ? _T_4006_24 : _T_5358_24; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_504 = _T_4557 ? _T_4006_25 : _T_5358_25; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_505 = _T_4557 ? _T_4006_26 : _T_5358_26; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_506 = _T_4557 ? _T_4006_27 : _T_5358_27; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_507 = _T_4557 ? _T_4006_28 : _T_5358_28; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_508 = _T_4557 ? _T_4006_29 : _T_5358_29; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_509 = _T_4557 ? _T_4006_30 : _T_5358_30; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_510 = _T_4557 ? _T_4006_31 : _T_5358_31; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_511 = _T_4557 ? _T_4006_32 : _T_5358_32; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_512 = _T_4557 ? _T_4006_33 : _T_5358_33; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_513 = _T_4557 ? _T_4006_34 : _T_5358_34; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_514 = _T_4557 ? _T_4006_35 : _T_5358_35; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_515 = _T_4557 ? _T_4006_36 : _T_5358_36; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_516 = _T_4557 ? _T_4006_37 : _T_5358_37; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_517 = _T_4557 ? _T_4006_38 : _T_5358_38; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_518 = _T_4557 ? _T_4006_39 : _T_5358_39; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_519 = _T_4557 ? _T_4006_40 : _T_5358_40; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_520 = _T_4557 ? _T_4006_41 : _T_5358_41; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_521 = _T_4557 ? _T_4006_42 : _T_5358_42; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_522 = _T_4557 ? _T_4006_43 : _T_5358_43; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_523 = _T_4557 ? _T_4006_44 : _T_5358_44; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_524 = _T_4557 ? _T_4006_45 : _T_5358_45; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_525 = _T_4557 ? _T_4006_46 : _T_5358_46; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_526 = _T_4557 ? _T_4006_47 : _T_5358_47; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_527 = _T_4557 ? _T_4006_48 : _T_5358_48; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_528 = _T_4557 ? _T_4006_49 : _T_5358_49; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_529 = _T_4557 ? _T_4006_50 : _T_5358_50; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_530 = _T_4557 ? _T_4006_51 : _T_5358_51; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_531 = _T_4557 ? _T_4006_52 : _T_5358_52; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_532 = _T_4557 ? _T_4006_53 : _T_5358_53; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_533 = _T_4557 ? _T_4006_54 : _T_5358_54; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_534 = _T_4557 ? _T_4006_55 : _T_5358_55; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_535 = _T_4557 ? _T_4006_56 : _T_5358_56; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_536 = _T_4557 ? _T_4006_57 : _T_5358_57; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_537 = _T_4557 ? _T_4006_58 : _T_5358_58; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_538 = _T_4557 ? _T_4006_59 : _T_5358_59; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_539 = _T_4557 ? _T_4006_60 : _T_5358_60; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_540 = _T_4557 ? _T_4006_61 : _T_5358_61; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_541 = _T_4557 ? _T_4006_62 : _T_5358_62; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_542 = _T_4557 ? _T_4006_63 : _T_5358_63; // @[Reg.scala 20:19:@3209.4]
  assign _T_5561 = {_T_5358_7,_T_5358_6,_T_5358_5,_T_5358_4,_T_5358_3,_T_5358_2,_T_5358_1,_T_5358_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3281.4]
  assign _T_5569 = {_T_5358_15,_T_5358_14,_T_5358_13,_T_5358_12,_T_5358_11,_T_5358_10,_T_5358_9,_T_5358_8,_T_5561}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3289.4]
  assign _T_5576 = {_T_5358_23,_T_5358_22,_T_5358_21,_T_5358_20,_T_5358_19,_T_5358_18,_T_5358_17,_T_5358_16}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3296.4]
  assign _T_5585 = {_T_5358_31,_T_5358_30,_T_5358_29,_T_5358_28,_T_5358_27,_T_5358_26,_T_5358_25,_T_5358_24,_T_5576,_T_5569}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3305.4]
  assign _T_5592 = {_T_5358_39,_T_5358_38,_T_5358_37,_T_5358_36,_T_5358_35,_T_5358_34,_T_5358_33,_T_5358_32}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3312.4]
  assign _T_5600 = {_T_5358_47,_T_5358_46,_T_5358_45,_T_5358_44,_T_5358_43,_T_5358_42,_T_5358_41,_T_5358_40,_T_5592}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3320.4]
  assign _T_5607 = {_T_5358_55,_T_5358_54,_T_5358_53,_T_5358_52,_T_5358_51,_T_5358_50,_T_5358_49,_T_5358_48}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3327.4]
  assign _T_5616 = {_T_5358_63,_T_5358_62,_T_5358_61,_T_5358_60,_T_5358_59,_T_5358_58,_T_5358_57,_T_5358_56,_T_5607,_T_5600}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3336.4]
  assign sc2cdma_dat_updt = _T_883; // @[NV_NVDLA_CSC_dl_for_check.scala 332:21:@326.4]
  assign sc2cdma_dat_entries = _T_889; // @[NV_NVDLA_CSC_dl_for_check.scala 334:24:@336.4]
  assign sc2cdma_dat_slices = _T_886; // @[NV_NVDLA_CSC_dl_for_check.scala 333:23:@331.4]
  assign sc2buf_dat_rd_en = _T_1495; // @[NV_NVDLA_CSC_dl_for_check.scala 749:29:@933.4]
  assign sc2buf_dat_rd_addr = _T_1502[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 750:28:@934.4]
  assign sc2mac_dat_a_valid = _T_4552; // @[NV_NVDLA_CSC_dl_for_check.scala 1198:23:@2929.4]
  assign sc2mac_dat_a_mask = {_T_5089,_T_5058}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:27:@3141.4]
  assign sc2mac_dat_a_data0 = _T_5619; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3343.4]
  assign sc2mac_dat_a_data1 = _T_5623; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3353.4]
  assign sc2mac_dat_a_data2 = _T_5627; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3363.4]
  assign sc2mac_dat_a_data3 = _T_5631; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3373.4]
  assign sc2mac_dat_a_data4 = _T_5635; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3383.4]
  assign sc2mac_dat_a_data5 = _T_5639; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3393.4]
  assign sc2mac_dat_a_data6 = _T_5643; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3403.4]
  assign sc2mac_dat_a_data7 = _T_5647; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3413.4]
  assign sc2mac_dat_a_data8 = _T_5651; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3423.4]
  assign sc2mac_dat_a_data9 = _T_5655; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3433.4]
  assign sc2mac_dat_a_data10 = _T_5659; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3443.4]
  assign sc2mac_dat_a_data11 = _T_5663; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3453.4]
  assign sc2mac_dat_a_data12 = _T_5667; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3463.4]
  assign sc2mac_dat_a_data13 = _T_5671; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3473.4]
  assign sc2mac_dat_a_data14 = _T_5675; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3483.4]
  assign sc2mac_dat_a_data15 = _T_5679; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3493.4]
  assign sc2mac_dat_a_data16 = _T_5683; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3503.4]
  assign sc2mac_dat_a_data17 = _T_5687; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3513.4]
  assign sc2mac_dat_a_data18 = _T_5691; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3523.4]
  assign sc2mac_dat_a_data19 = _T_5695; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3533.4]
  assign sc2mac_dat_a_data20 = _T_5699; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3543.4]
  assign sc2mac_dat_a_data21 = _T_5703; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3553.4]
  assign sc2mac_dat_a_data22 = _T_5707; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3563.4]
  assign sc2mac_dat_a_data23 = _T_5711; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3573.4]
  assign sc2mac_dat_a_data24 = _T_5715; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3583.4]
  assign sc2mac_dat_a_data25 = _T_5719; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3593.4]
  assign sc2mac_dat_a_data26 = _T_5723; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3603.4]
  assign sc2mac_dat_a_data27 = _T_5727; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3613.4]
  assign sc2mac_dat_a_data28 = _T_5731; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3623.4]
  assign sc2mac_dat_a_data29 = _T_5735; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3633.4]
  assign sc2mac_dat_a_data30 = _T_5739; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3643.4]
  assign sc2mac_dat_a_data31 = _T_5743; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3653.4]
  assign sc2mac_dat_a_data32 = _T_5747; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3663.4]
  assign sc2mac_dat_a_data33 = _T_5751; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3673.4]
  assign sc2mac_dat_a_data34 = _T_5755; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3683.4]
  assign sc2mac_dat_a_data35 = _T_5759; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3693.4]
  assign sc2mac_dat_a_data36 = _T_5763; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3703.4]
  assign sc2mac_dat_a_data37 = _T_5767; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3713.4]
  assign sc2mac_dat_a_data38 = _T_5771; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3723.4]
  assign sc2mac_dat_a_data39 = _T_5775; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3733.4]
  assign sc2mac_dat_a_data40 = _T_5779; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3743.4]
  assign sc2mac_dat_a_data41 = _T_5783; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3753.4]
  assign sc2mac_dat_a_data42 = _T_5787; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3763.4]
  assign sc2mac_dat_a_data43 = _T_5791; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3773.4]
  assign sc2mac_dat_a_data44 = _T_5795; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3783.4]
  assign sc2mac_dat_a_data45 = _T_5799; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3793.4]
  assign sc2mac_dat_a_data46 = _T_5803; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3803.4]
  assign sc2mac_dat_a_data47 = _T_5807; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3813.4]
  assign sc2mac_dat_a_data48 = _T_5811; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3823.4]
  assign sc2mac_dat_a_data49 = _T_5815; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3833.4]
  assign sc2mac_dat_a_data50 = _T_5819; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3843.4]
  assign sc2mac_dat_a_data51 = _T_5823; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3853.4]
  assign sc2mac_dat_a_data52 = _T_5827; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3863.4]
  assign sc2mac_dat_a_data53 = _T_5831; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3873.4]
  assign sc2mac_dat_a_data54 = _T_5835; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3883.4]
  assign sc2mac_dat_a_data55 = _T_5839; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3893.4]
  assign sc2mac_dat_a_data56 = _T_5843; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3903.4]
  assign sc2mac_dat_a_data57 = _T_5847; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3913.4]
  assign sc2mac_dat_a_data58 = _T_5851; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3923.4]
  assign sc2mac_dat_a_data59 = _T_5855; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3933.4]
  assign sc2mac_dat_a_data60 = _T_5859; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3943.4]
  assign sc2mac_dat_a_data61 = _T_5863; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3953.4]
  assign sc2mac_dat_a_data62 = _T_5867; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3963.4]
  assign sc2mac_dat_a_data63 = _T_5871; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3973.4]
  assign sc2mac_dat_a_pd = _T_4559; // @[NV_NVDLA_CSC_dl_for_check.scala 1200:25:@2938.4]
  assign sc2mac_dat_b_valid = _T_4555; // @[NV_NVDLA_CSC_dl_for_check.scala 1199:23:@2932.4]
  assign sc2mac_dat_b_mask = {_T_5616,_T_5585}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:27:@3338.4]
  assign sc2mac_dat_b_data0 = _T_5621; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3348.4]
  assign sc2mac_dat_b_data1 = _T_5625; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3358.4]
  assign sc2mac_dat_b_data2 = _T_5629; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3368.4]
  assign sc2mac_dat_b_data3 = _T_5633; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3378.4]
  assign sc2mac_dat_b_data4 = _T_5637; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3388.4]
  assign sc2mac_dat_b_data5 = _T_5641; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3398.4]
  assign sc2mac_dat_b_data6 = _T_5645; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3408.4]
  assign sc2mac_dat_b_data7 = _T_5649; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3418.4]
  assign sc2mac_dat_b_data8 = _T_5653; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3428.4]
  assign sc2mac_dat_b_data9 = _T_5657; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3438.4]
  assign sc2mac_dat_b_data10 = _T_5661; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3448.4]
  assign sc2mac_dat_b_data11 = _T_5665; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3458.4]
  assign sc2mac_dat_b_data12 = _T_5669; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3468.4]
  assign sc2mac_dat_b_data13 = _T_5673; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3478.4]
  assign sc2mac_dat_b_data14 = _T_5677; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3488.4]
  assign sc2mac_dat_b_data15 = _T_5681; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3498.4]
  assign sc2mac_dat_b_data16 = _T_5685; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3508.4]
  assign sc2mac_dat_b_data17 = _T_5689; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3518.4]
  assign sc2mac_dat_b_data18 = _T_5693; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3528.4]
  assign sc2mac_dat_b_data19 = _T_5697; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3538.4]
  assign sc2mac_dat_b_data20 = _T_5701; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3548.4]
  assign sc2mac_dat_b_data21 = _T_5705; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3558.4]
  assign sc2mac_dat_b_data22 = _T_5709; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3568.4]
  assign sc2mac_dat_b_data23 = _T_5713; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3578.4]
  assign sc2mac_dat_b_data24 = _T_5717; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3588.4]
  assign sc2mac_dat_b_data25 = _T_5721; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3598.4]
  assign sc2mac_dat_b_data26 = _T_5725; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3608.4]
  assign sc2mac_dat_b_data27 = _T_5729; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3618.4]
  assign sc2mac_dat_b_data28 = _T_5733; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3628.4]
  assign sc2mac_dat_b_data29 = _T_5737; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3638.4]
  assign sc2mac_dat_b_data30 = _T_5741; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3648.4]
  assign sc2mac_dat_b_data31 = _T_5745; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3658.4]
  assign sc2mac_dat_b_data32 = _T_5749; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3668.4]
  assign sc2mac_dat_b_data33 = _T_5753; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3678.4]
  assign sc2mac_dat_b_data34 = _T_5757; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3688.4]
  assign sc2mac_dat_b_data35 = _T_5761; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3698.4]
  assign sc2mac_dat_b_data36 = _T_5765; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3708.4]
  assign sc2mac_dat_b_data37 = _T_5769; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3718.4]
  assign sc2mac_dat_b_data38 = _T_5773; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3728.4]
  assign sc2mac_dat_b_data39 = _T_5777; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3738.4]
  assign sc2mac_dat_b_data40 = _T_5781; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3748.4]
  assign sc2mac_dat_b_data41 = _T_5785; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3758.4]
  assign sc2mac_dat_b_data42 = _T_5789; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3768.4]
  assign sc2mac_dat_b_data43 = _T_5793; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3778.4]
  assign sc2mac_dat_b_data44 = _T_5797; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3788.4]
  assign sc2mac_dat_b_data45 = _T_5801; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3798.4]
  assign sc2mac_dat_b_data46 = _T_5805; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3808.4]
  assign sc2mac_dat_b_data47 = _T_5809; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3818.4]
  assign sc2mac_dat_b_data48 = _T_5813; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3828.4]
  assign sc2mac_dat_b_data49 = _T_5817; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3838.4]
  assign sc2mac_dat_b_data50 = _T_5821; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3848.4]
  assign sc2mac_dat_b_data51 = _T_5825; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3858.4]
  assign sc2mac_dat_b_data52 = _T_5829; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3868.4]
  assign sc2mac_dat_b_data53 = _T_5833; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3878.4]
  assign sc2mac_dat_b_data54 = _T_5837; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3888.4]
  assign sc2mac_dat_b_data55 = _T_5841; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3898.4]
  assign sc2mac_dat_b_data56 = _T_5845; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3908.4]
  assign sc2mac_dat_b_data57 = _T_5849; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3918.4]
  assign sc2mac_dat_b_data58 = _T_5853; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3928.4]
  assign sc2mac_dat_b_data59 = _T_5857; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3938.4]
  assign sc2mac_dat_b_data60 = _T_5861; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3948.4]
  assign sc2mac_dat_b_data61 = _T_5865; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3958.4]
  assign sc2mac_dat_b_data62 = _T_5869; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3968.4]
  assign sc2mac_dat_b_data63 = _T_5873; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3978.4]
  assign sc2mac_dat_b_pd = _T_4563; // @[NV_NVDLA_CSC_dl_for_check.scala 1201:25:@2944.4]
  assign slcg_wg_en = 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 273:15:@243.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_432 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_439 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_446 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_453 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_460 = _RAND_4[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_467 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_474 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_488 = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_495 = _RAND_8[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_502 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_509 = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_548 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_555 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_562 = _RAND_13[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_569 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_576 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_583 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_586 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_589 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_595 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_598 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_601 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_604 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_610 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_613 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_619 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_622 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_625 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_632 = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_639 = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_649 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_656 = _RAND_31[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_663 = _RAND_32[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_670 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_677 = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_684 = _RAND_35[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_691 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_698 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_705 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_712 = _RAND_39[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_719 = _RAND_40[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_726 = _RAND_41[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_733 = _RAND_42[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_740 = _RAND_43[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_793 = _RAND_44[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_1934 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_1928 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_1925 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1948 = _RAND_48[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1942 = _RAND_49[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1939 = _RAND_50[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_883 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_886 = _RAND_52[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_889 = _RAND_53[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_894 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_897 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_900 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_903 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_906 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_928 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_931 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_934 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_937 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_942 = _RAND_63[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_945 = _RAND_64[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_948 = _RAND_65[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_951 = _RAND_66[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_996 = _RAND_67[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1007 = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1023 = _RAND_69[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1052 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1046 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1049 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1078 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1083 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1086 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1107 = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1121 = _RAND_77[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1124 = _RAND_78[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1127 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1130 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1133 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1136 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1141 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1144 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1256 = _RAND_85[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1259 = _RAND_86[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1333 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1336 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1339 = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1342 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1345 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1348 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1351 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1354 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1357 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1360 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1365 = _RAND_97[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1368 = _RAND_98[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1371 = _RAND_99[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1374 = _RAND_100[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1377 = _RAND_101[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1380 = _RAND_102[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1383 = _RAND_103[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1476_0 = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1476_1 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1476_2 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1476_3 = _RAND_107[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1495 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1502 = _RAND_109[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1505 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1511 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1514 = _RAND_112[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1517 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1520 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1523 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_1526 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_1529 = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_1532 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_1535 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1538 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1660 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1663 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1666 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1669 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_1672 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1675 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1680 = _RAND_127[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1683 = _RAND_128[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1686 = _RAND_129[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1689 = _RAND_130[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1692 = _RAND_131[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1695 = _RAND_132[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_1768 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_1780 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {16{`RANDOM}};
  _T_1791 = _RAND_135[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {16{`RANDOM}};
  _T_1799 = _RAND_136[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_1899 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_1902 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_1905 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_1908 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_1911 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_1914 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_1917 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_1920 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_1931 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_1945 = _RAND_146[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {8{`RANDOM}};
  _T_2328 = _RAND_147[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {4{`RANDOM}};
  _T_2330 = _RAND_148[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {4{`RANDOM}};
  _T_2332 = _RAND_149[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {4{`RANDOM}};
  _T_2334 = _RAND_150[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {4{`RANDOM}};
  _T_2336 = _RAND_151[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {4{`RANDOM}};
  _T_2338 = _RAND_152[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_3136 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_3406_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_3406_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_3406_2 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_3406_3 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_3406_4 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_3406_5 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_3406_6 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_3406_7 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_3406_8 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_3406_9 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_3406_10 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_3406_11 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_3406_12 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_3406_13 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_3406_14 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_3406_15 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_3406_16 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_3406_17 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_3406_18 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_3406_19 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_3406_20 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_3406_21 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_3406_22 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_3406_23 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_3406_24 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_3406_25 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_3406_26 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_3406_27 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_3406_28 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_3406_29 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_3406_30 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_3406_31 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_3406_32 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_3406_33 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_3406_34 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_3406_35 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_3406_36 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_3406_37 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_3406_38 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_3406_39 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_3406_40 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_3406_41 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_3406_42 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_3406_43 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_3406_44 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_3406_45 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_3406_46 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_3406_47 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_3406_48 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_3406_49 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_3406_50 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_3406_51 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_3406_52 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_3406_53 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_3406_54 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_3406_55 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_3406_56 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_3406_57 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_3406_58 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_3406_59 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_3406_60 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_3406_61 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_3406_62 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_3406_63 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_3606_0 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_3606_1 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_3606_2 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_3606_3 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_3606_4 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_3606_5 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_3606_6 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_3606_7 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_3606_8 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_3606_9 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_3606_10 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3606_11 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3606_12 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3606_13 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3606_14 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3606_15 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3606_16 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3606_17 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3606_18 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3606_19 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3606_20 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3606_21 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3606_22 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3606_23 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3606_24 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3606_25 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3606_26 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3606_27 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3606_28 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3606_29 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3606_30 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3606_31 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3606_32 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3606_33 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3606_34 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3606_35 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3606_36 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3606_37 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3606_38 = _RAND_256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3606_39 = _RAND_257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_3606_40 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_3606_41 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_3606_42 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_3606_43 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_3606_44 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_3606_45 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_3606_46 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_3606_47 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_3606_48 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_3606_49 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_3606_50 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_3606_51 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_3606_52 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_3606_53 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_3606_54 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_3606_55 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_3606_56 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_3606_57 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_3606_58 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_3606_59 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_3606_60 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_3606_61 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_3606_62 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_3606_63 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_3739 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_4006_0 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_4006_1 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_4006_2 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_4006_3 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_4006_4 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_4006_5 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_4006_6 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_4006_7 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_4006_8 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_4006_9 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_4006_10 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_4006_11 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_4006_12 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_4006_13 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_4006_14 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_4006_15 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_4006_16 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_4006_17 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_4006_18 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_4006_19 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_4006_20 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_4006_21 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_4006_22 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_4006_23 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_4006_24 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_4006_25 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_4006_26 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_4006_27 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_4006_28 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_4006_29 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_4006_30 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_4006_31 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_4006_32 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_4006_33 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_4006_34 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_4006_35 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_4006_36 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_4006_37 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_4006_38 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_4006_39 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_4006_40 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_4006_41 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_4006_42 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_4006_43 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_4006_44 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_4006_45 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_4006_46 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_4006_47 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_4006_48 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_4006_49 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_4006_50 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_4006_51 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_4006_52 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_4006_53 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_4006_54 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_4006_55 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_4006_56 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_4006_57 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_4006_58 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_4006_59 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_4006_60 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_4006_61 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_4006_62 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_4006_63 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_4205 = _RAND_347[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_4209_0 = _RAND_348[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_4209_1 = _RAND_349[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_4209_2 = _RAND_350[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_4209_3 = _RAND_351[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_4209_4 = _RAND_352[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_4209_5 = _RAND_353[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_4209_6 = _RAND_354[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_4209_7 = _RAND_355[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_4209_8 = _RAND_356[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_4209_9 = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_4209_10 = _RAND_358[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4209_11 = _RAND_359[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4209_12 = _RAND_360[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4209_13 = _RAND_361[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4209_14 = _RAND_362[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4209_15 = _RAND_363[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4209_16 = _RAND_364[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4209_17 = _RAND_365[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4209_18 = _RAND_366[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4209_19 = _RAND_367[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4209_20 = _RAND_368[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4209_21 = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4209_22 = _RAND_370[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4209_23 = _RAND_371[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4209_24 = _RAND_372[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4209_25 = _RAND_373[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4209_26 = _RAND_374[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4209_27 = _RAND_375[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4209_28 = _RAND_376[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4209_29 = _RAND_377[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4209_30 = _RAND_378[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4209_31 = _RAND_379[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4209_32 = _RAND_380[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4209_33 = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4209_34 = _RAND_382[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4209_35 = _RAND_383[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4209_36 = _RAND_384[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4209_37 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4209_38 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4209_39 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4209_40 = _RAND_388[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4209_41 = _RAND_389[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4209_42 = _RAND_390[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4209_43 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4209_44 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4209_45 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4209_46 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4209_47 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4209_48 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4209_49 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4209_50 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4209_51 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4209_52 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4209_53 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4209_54 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4209_55 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4209_56 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4209_57 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4209_58 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4209_59 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4209_60 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4209_61 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4209_62 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4209_63 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4546 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4552 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4555 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4559 = _RAND_415[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4563 = _RAND_416[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_4831_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_4831_1 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_4831_2 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_4831_3 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_4831_4 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_4831_5 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_4831_6 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_4831_7 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_4831_8 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_4831_9 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_4831_10 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_4831_11 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_4831_12 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_4831_13 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_4831_14 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_4831_15 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_4831_16 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_4831_17 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_4831_18 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_4831_19 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_4831_20 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_4831_21 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_4831_22 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_4831_23 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_4831_24 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_4831_25 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_4831_26 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_4831_27 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_4831_28 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_4831_29 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_4831_30 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_4831_31 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_4831_32 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_4831_33 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_4831_34 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_4831_35 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_4831_36 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_4831_37 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_4831_38 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_4831_39 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_4831_40 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_4831_41 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_4831_42 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_4831_43 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_4831_44 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_4831_45 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_4831_46 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_4831_47 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_4831_48 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_4831_49 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_4831_50 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_4831_51 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_4831_52 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_4831_53 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_4831_54 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_4831_55 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_4831_56 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_4831_57 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_4831_58 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_4831_59 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_4831_60 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_4831_61 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_4831_62 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_4831_63 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_5358_0 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_5358_1 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_5358_2 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_5358_3 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_5358_4 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_5358_5 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_5358_6 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_5358_7 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_5358_8 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_5358_9 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_5358_10 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_5358_11 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_5358_12 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_5358_13 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_5358_14 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_5358_15 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_5358_16 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_5358_17 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_5358_18 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_5358_19 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_5358_20 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_5358_21 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_5358_22 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_5358_23 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_5358_24 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_5358_25 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_5358_26 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_5358_27 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_5358_28 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_5358_29 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_5358_30 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_5358_31 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_5358_32 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_5358_33 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_5358_34 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_5358_35 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_5358_36 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_5358_37 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_5358_38 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_5358_39 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_5358_40 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_5358_41 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_5358_42 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_5358_43 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_5358_44 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_5358_45 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_5358_46 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_5358_47 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_5358_48 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_5358_49 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_5358_50 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_5358_51 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_5358_52 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_5358_53 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_5358_54 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_5358_55 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_5358_56 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_5358_57 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_5358_58 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_5358_59 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_5358_60 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_5358_61 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_5358_62 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_5358_63 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5619 = _RAND_545[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5621 = _RAND_546[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5623 = _RAND_547[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5625 = _RAND_548[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5627 = _RAND_549[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_5629 = _RAND_550[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_5631 = _RAND_551[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_5633 = _RAND_552[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_5635 = _RAND_553[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_5637 = _RAND_554[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_5639 = _RAND_555[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_5641 = _RAND_556[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_5643 = _RAND_557[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_5645 = _RAND_558[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_5647 = _RAND_559[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_5649 = _RAND_560[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_5651 = _RAND_561[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_5653 = _RAND_562[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_5655 = _RAND_563[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_5657 = _RAND_564[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_5659 = _RAND_565[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_5661 = _RAND_566[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_5663 = _RAND_567[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_5665 = _RAND_568[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_5667 = _RAND_569[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_5669 = _RAND_570[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_5671 = _RAND_571[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_5673 = _RAND_572[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_5675 = _RAND_573[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_5677 = _RAND_574[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_5679 = _RAND_575[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_5681 = _RAND_576[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_5683 = _RAND_577[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_5685 = _RAND_578[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_5687 = _RAND_579[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_5689 = _RAND_580[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_5691 = _RAND_581[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_5693 = _RAND_582[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_5695 = _RAND_583[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_5697 = _RAND_584[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_5699 = _RAND_585[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_5701 = _RAND_586[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_5703 = _RAND_587[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_5705 = _RAND_588[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_5707 = _RAND_589[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_5709 = _RAND_590[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_5711 = _RAND_591[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_5713 = _RAND_592[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_5715 = _RAND_593[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_5717 = _RAND_594[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_5719 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_5721 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_5723 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_5725 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_5727 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_5729 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_5731 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_5733 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_5735 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_5737 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_5739 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_5741 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_5743 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_5745 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_5747 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_5749 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_5751 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_5753 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_5755 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_5757 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_5759 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_5761 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_5763 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_5765 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_5767 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_5769 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_5771 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_5773 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_5775 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_5777 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_5779 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_5781 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_5783 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_5785 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_5787 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_5789 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_5791 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_5793 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_5795 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_5797 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_5799 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_5801 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_5803 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_5805 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_5807 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_5809 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_5811 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_5813 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_5815 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_5817 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_5819 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_5821 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_5823 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_5825 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_5827 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_5829 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_5831 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_5833 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_5835 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_5837 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_5839 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_5841 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_5843 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_5845 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_5847 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_5849 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_5851 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_5853 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_5855 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_5857 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_5859 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_5861 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_5863 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_5865 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_5867 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_5869 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_5871 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_5873 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge nvdla_core_clk) begin
    if (_T_337) begin
      _T_432 <= 1'h0;
    end else begin
      _T_432 <= _T_347;
    end
    if (_T_337) begin
      _T_439 <= 6'h0;
    end else begin
      if (_T_347) begin
        _T_439 <= 6'h1;
      end
    end
    if (_T_337) begin
      _T_446 <= 14'h0;
    end else begin
      if (_T_347) begin
        _T_446 <= {{2'd0}, _T_522};
      end
    end
    if (_T_337) begin
      _T_453 <= 14'h0;
    end else begin
      if (_T_347) begin
        _T_453 <= {{2'd0}, _T_515};
      end
    end
    if (_T_337) begin
      _T_460 <= 15'h0;
    end else begin
      if (_T_347) begin
        _T_460 <= _T_511;
      end
    end
    if (_T_337) begin
      _T_467 <= 15'h0;
    end else begin
      if (_T_347) begin
        _T_467 <= _T_514;
      end
    end
    if (_T_337) begin
      _T_474 <= 13'h0;
    end else begin
      if (_T_347) begin
        _T_474 <= reg2dp_dataout_width;
      end
    end
    if (_T_337) begin
      _T_488 <= 15'h0;
    end else begin
      if (_T_432) begin
        _T_488 <= _T_530;
      end
    end
    if (_T_337) begin
      _T_495 <= 12'h0;
    end else begin
      if (_T_432) begin
        _T_495 <= _T_517;
      end
    end
    if (_T_337) begin
      _T_502 <= 12'h0;
    end else begin
      if (_T_432) begin
        _T_502 <= _T_519;
      end
    end
    if (_T_337) begin
      _T_509 <= 14'h0;
    end else begin
      if (_T_347) begin
        if (reg2dp_skip_data_rls) begin
          _T_509 <= _T_524;
        end else begin
          _T_509 <= _T_526;
        end
      end
    end
    if (_T_337) begin
      _T_548 <= 34'h0;
    end else begin
      if (_T_347) begin
        if (_T_352) begin
          _T_548 <= 34'h3ffffffff;
        end else begin
          _T_548 <= 34'h0;
        end
      end
    end
    if (_T_337) begin
      _T_555 <= 5'h0;
    end else begin
      if (_T_347) begin
        _T_555 <= _T_758;
      end
    end
    if (_T_337) begin
      _T_562 <= 14'h0;
    end else begin
      if (_T_347) begin
        _T_562 <= _T_760;
      end
    end
    if (_T_337) begin
      _T_569 <= 13'h0;
    end else begin
      if (_T_347) begin
        _T_569 <= reg2dp_datain_width_ext;
      end
    end
    if (_T_337) begin
      _T_576 <= 13'h0;
    end else begin
      if (_T_347) begin
        _T_576 <= reg2dp_datain_height_ext;
      end
    end
    if (_T_337) begin
      _T_583 <= 11'h0;
    end else begin
      if (_T_347) begin
        _T_583 <= _T_767;
      end
    end
    if (_T_337) begin
      _T_586 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_586 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_589 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_589 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_595 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_595 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_598 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_598 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_601 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_601 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_604 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_604 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_610 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_610 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_613 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_613 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_619 <= 3'h1;
    end else begin
      if (_T_347) begin
        _T_619 <= _T_360;
      end
    end
    if (_T_337) begin
      _T_622 <= 3'h1;
    end else begin
      if (_T_347) begin
        if (_T_352) begin
          _T_622 <= _T_360;
        end else begin
          _T_622 <= 3'h1;
        end
      end
    end
    if (_T_337) begin
      _T_625 <= 3'h1;
    end else begin
      if (_T_347) begin
        if (_T_352) begin
          _T_625 <= _T_360;
        end else begin
          _T_625 <= 3'h1;
        end
      end
    end
    if (_T_337) begin
      _T_632 <= 4'h0;
    end else begin
      if (_T_347) begin
        _T_632 <= _T_367;
      end
    end
    if (_T_337) begin
      _T_639 <= 4'h0;
    end else begin
      if (_T_347) begin
        _T_639 <= _T_421;
      end
    end
    if (_T_337) begin
      _T_649 <= 5'h0;
    end else begin
      if (_T_347) begin
        _T_649 <= 5'h0;
      end
    end
    if (_T_337) begin
      _T_656 <= 7'h0;
    end else begin
      if (_T_347) begin
        if (_T_403) begin
          _T_656 <= _T_396;
        end else begin
          _T_656 <= {{1'd0}, _T_402};
        end
      end
    end
    if (_T_337) begin
      _T_663 <= 7'h0;
    end else begin
      if (_T_347) begin
        _T_663 <= _T_407;
      end
    end
    if (_T_337) begin
      _T_670 <= 8'h0;
    end else begin
      if (_T_347) begin
        if (_T_403) begin
          _T_670 <= _T_410;
        end else begin
          _T_670 <= {{1'd0}, _T_415};
        end
      end
    end
    if (_T_337) begin
      _T_677 <= 7'h0;
    end else begin
      if (_T_347) begin
        _T_677 <= {{1'd0}, _T_379};
      end
    end
    if (_T_337) begin
      _T_684 <= 12'h0;
    end else begin
      if (_T_347) begin
        _T_684 <= _T_419;
      end
    end
    if (_T_337) begin
      _T_691 <= 6'h0;
    end else begin
      if (_T_347) begin
        if (_T_352) begin
          _T_691 <= 6'h1;
        end else begin
          _T_691 <= _T_424;
        end
      end
    end
    if (_T_337) begin
      _T_698 <= 6'h0;
    end else begin
      if (_T_347) begin
        if (_T_352) begin
          _T_698 <= 6'h1;
        end else begin
          _T_698 <= _T_428;
        end
      end
    end
    if (_T_337) begin
      _T_705 <= 16'h0;
    end else begin
      if (_T_347) begin
        _T_705 <= reg2dp_pad_value;
      end
    end
    if (_T_337) begin
      _T_712 <= 15'h0;
    end else begin
      if (_T_347) begin
        _T_712 <= _T_771;
      end
    end
    if (_T_337) begin
      _T_719 <= 15'h0;
    end else begin
      if (_T_432) begin
        _T_719 <= _T_460;
      end
    end
    if (_T_337) begin
      _T_726 <= 15'h0;
    end else begin
      if (_T_432) begin
        _T_726 <= _T_460;
      end
    end
    if (_T_337) begin
      _T_733 <= 14'h0;
    end else begin
      if (_T_343) begin
        _T_733 <= _T_509;
      end
    end
    if (_T_337) begin
      _T_740 <= 15'h0;
    end else begin
      if (_T_343) begin
        _T_740 <= _T_530;
      end
    end
    if (_T_337) begin
      _T_1934 <= 1'h0;
    end else begin
      _T_1934 <= _T_1931;
    end
    if (_T_337) begin
      _T_1928 <= 1'h0;
    end else begin
      _T_1928 <= _T_1925;
    end
    if (_T_337) begin
      _T_1925 <= 1'h0;
    end else begin
      _T_1925 <= _T_1675;
    end
    if (_T_337) begin
      _T_1948 <= 27'h0;
    end else begin
      if (_T_1931) begin
        _T_1948 <= _T_1945;
      end
    end
    if (_T_337) begin
      _T_1942 <= 27'h0;
    end else begin
      if (_T_1925) begin
        _T_1942 <= _T_1939;
      end
    end
    if (_T_337) begin
      _T_1939 <= 27'h0;
    end else begin
      if (_T_1675) begin
        _T_1939 <= _T_1957;
      end
    end
    if (_T_337) begin
      _T_883 <= 1'h0;
    end else begin
      _T_883 <= _T_878;
    end
    if (_T_337) begin
      _T_886 <= 14'h0;
    end else begin
      if (_T_878) begin
        if (_T_871) begin
          _T_886 <= _T_446;
        end else begin
          _T_886 <= _T_733;
        end
      end
    end
    if (_T_337) begin
      _T_889 <= 15'h0;
    end else begin
      if (_T_878) begin
        if (_T_871) begin
          _T_889 <= _T_488;
        end else begin
          _T_889 <= _T_740;
        end
      end
    end
    if (_T_337) begin
      _T_894 <= 1'h0;
    end else begin
      _T_894 <= sg2dl_pvld;
    end
    if (_T_337) begin
      _T_897 <= 1'h0;
    end else begin
      _T_897 <= _T_894;
    end
    if (_T_337) begin
      _T_900 <= 1'h0;
    end else begin
      _T_900 <= _T_897;
    end
    if (_T_337) begin
      _T_903 <= 1'h0;
    end else begin
      _T_903 <= _T_900;
    end
    if (_T_337) begin
      _T_906 <= 1'h0;
    end else begin
      _T_906 <= _T_903;
    end
    if (_T_337) begin
      _T_928 <= 1'h0;
    end else begin
      _T_928 <= _T_906;
    end
    if (_T_337) begin
      _T_931 <= 1'h0;
    end else begin
      _T_931 <= _T_928;
    end
    if (_T_337) begin
      _T_934 <= 1'h0;
    end else begin
      _T_934 <= _T_931;
    end
    if (_T_337) begin
      _T_937 <= 1'h0;
    end else begin
      _T_937 <= _T_934;
    end
    if (_T_337) begin
      _T_942 <= 31'h0;
    end else begin
      if (_T_906) begin
        _T_942 <= _T_939;
      end
    end
    if (_T_337) begin
      _T_945 <= 31'h0;
    end else begin
      if (_T_928) begin
        _T_945 <= _T_942;
      end
    end
    if (_T_337) begin
      _T_948 <= 31'h0;
    end else begin
      if (_T_931) begin
        _T_948 <= _T_945;
      end
    end
    if (_T_337) begin
      _T_951 <= 31'h0;
    end else begin
      if (_T_934) begin
        _T_951 <= _T_948;
      end
    end
    if (_T_337) begin
      _T_996 <= 5'h0;
    end else begin
      if (_T_347) begin
        _T_996 <= 5'h0;
      end else begin
        if (_T_1004) begin
          _T_996 <= 5'h0;
        end else begin
          _T_996 <= _T_1001;
        end
      end
    end
    if (_T_337) begin
      _T_1007 <= 2'h0;
    end else begin
      if (_T_1017) begin
        if (_T_1018) begin
          _T_1007 <= 2'h0;
        end else begin
          _T_1007 <= _T_1012;
        end
      end
    end
    if (_T_337) begin
      _T_1023 <= 7'h0;
    end else begin
      if (_T_1035) begin
        if (_T_347) begin
          _T_1023 <= 7'h0;
        end else begin
          if (_T_1038) begin
            _T_1023 <= 7'h0;
          end else begin
            if (_T_1033) begin
              _T_1023 <= 7'h0;
            end else begin
              _T_1023 <= _T_1030;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1052 <= 1'h0;
    end else begin
      if (_T_959) begin
        _T_1052 <= 1'h1;
      end else begin
        if (_T_1072) begin
          _T_1052 <= 1'h0;
        end
      end
    end
    if (_T_337) begin
      _T_1046 <= 1'h0;
    end else begin
      if (_T_1055) begin
        _T_1046 <= 1'h0;
      end else begin
        if (_T_959) begin
          _T_1046 <= 1'h1;
        end
      end
    end
    if (_T_337) begin
      _T_1049 <= 1'h0;
    end else begin
      _T_1049 <= _T_1060;
    end
    if (_T_337) begin
      _T_1078 <= 8'h0;
    end else begin
      if (_T_1075) begin
        _T_1078 <= _T_1080;
      end
    end
    if (_T_337) begin
      _T_1083 <= 13'h0;
    end else begin
      if (_T_1101) begin
        if (_T_347) begin
          _T_1083 <= {{9'd0}, _T_365};
        end else begin
          if (_T_1095) begin
            _T_1083 <= _T_1086;
          end else begin
            if (_T_1091) begin
              _T_1083 <= {{9'd0}, _T_365};
            end else begin
              _T_1083 <= _T_1088;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1086 <= 13'h0;
    end else begin
      if (_T_1104) begin
        if (_T_347) begin
          _T_1086 <= {{9'd0}, _T_365};
        end else begin
          if (!(_T_1095)) begin
            if (_T_1091) begin
              _T_1086 <= {{9'd0}, _T_365};
            end else begin
              _T_1086 <= _T_1088;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1107 <= 11'h0;
    end else begin
      if (_T_1111) begin
        if (_T_347) begin
          _T_1107 <= 11'h0;
        end else begin
          if (_T_986) begin
            _T_1107 <= 11'h0;
          end else begin
            _T_1107 <= _T_1116;
          end
        end
      end
    end
    if (_T_337) begin
      _T_1121 <= 14'h0;
    end else begin
      if (_T_1165) begin
        if (_T_347) begin
          if (_T_352) begin
            _T_1121 <= 14'h0;
          end else begin
            _T_1121 <= _T_1148;
          end
        end else begin
          if (_T_1095) begin
            _T_1121 <= _T_1124;
          end else begin
            if (_T_1091) begin
              if (_T_352) begin
                _T_1121 <= 14'h0;
              end else begin
                _T_1121 <= _T_1148;
              end
            end else begin
              _T_1121 <= _T_1151;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1124 <= 14'h0;
    end else begin
      if (_T_1171) begin
        if (_T_347) begin
          if (_T_352) begin
            _T_1124 <= 14'h0;
          end else begin
            _T_1124 <= _T_1148;
          end
        end else begin
          if (!(_T_1095)) begin
            if (_T_1091) begin
              if (_T_352) begin
                _T_1124 <= 14'h0;
              end else begin
                _T_1124 <= _T_1148;
              end
            end else begin
              _T_1124 <= _T_1151;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1127 <= 16'h0;
    end else begin
      if (_T_1165) begin
        if (_T_432) begin
          _T_1127 <= {{9'd0}, _T_656};
        end else begin
          if (_T_1194) begin
            _T_1127 <= {{9'd0}, _T_656};
          end else begin
            if (_T_1198) begin
              _T_1127 <= _T_1200;
            end else begin
              if (_T_1202) begin
                _T_1127 <= _T_1204;
              end else begin
                if (_T_1207) begin
                  _T_1127 <= _T_1210;
                end else begin
                  if (_T_1212) begin
                    _T_1127 <= _T_1130;
                  end else begin
                    _T_1127 <= _T_1214;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1130 <= 16'h0;
    end else begin
      if (_T_1171) begin
        if (_T_432) begin
          _T_1130 <= {{9'd0}, _T_656};
        end else begin
          if (_T_1194) begin
            _T_1130 <= {{9'd0}, _T_656};
          end else begin
            if (_T_1198) begin
              _T_1130 <= _T_1200;
            end else begin
              if (_T_1202) begin
                _T_1130 <= _T_1204;
              end else begin
                if (_T_1207) begin
                  _T_1130 <= _T_1210;
                end else begin
                  if (!(_T_1212)) begin
                    _T_1130 <= _T_1214;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1133 <= 16'h0;
    end else begin
      if (_T_1243) begin
        if (_T_432) begin
          _T_1133 <= {{9'd0}, _T_656};
        end else begin
          if (_T_1194) begin
            _T_1133 <= {{9'd0}, _T_656};
          end else begin
            if (_T_1198) begin
              _T_1133 <= _T_1200;
            end else begin
              if (_T_1202) begin
                _T_1133 <= _T_1204;
              end else begin
                if (_T_1207) begin
                  _T_1133 <= _T_1210;
                end else begin
                  if (_T_1212) begin
                    _T_1133 <= _T_1130;
                  end else begin
                    _T_1133 <= _T_1214;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1136 <= 13'h2;
    end else begin
      if (_T_1183) begin
        _T_1136 <= 13'h2;
      end else begin
        if (_T_1185) begin
          _T_1136 <= _T_1188;
        end
      end
    end
    if (_T_337) begin
      _T_1141 <= 1'h0;
    end else begin
      if (_T_1075) begin
        _T_1141 <= _T_1253;
      end
    end
    if (_T_337) begin
      _T_1144 <= 1'h0;
    end else begin
      if (_T_1075) begin
        if (_T_1245) begin
          _T_1144 <= 1'h1;
        end else begin
          if (_T_1141) begin
            _T_1144 <= 1'h0;
          end
        end
      end
    end
    if (_T_337) begin
      _T_1256 <= 14'h0;
    end else begin
      if (_T_1277) begin
        if (_T_1267) begin
          _T_1256 <= _T_1263;
        end else begin
          if (_T_1095) begin
            _T_1256 <= _T_1259;
          end else begin
            if (_T_1091) begin
              _T_1256 <= _T_1265;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1259 <= 14'h0;
    end else begin
      if (_T_1104) begin
        if (_T_1267) begin
          _T_1259 <= _T_1263;
        end else begin
          if (!(_T_1095)) begin
            if (_T_1091) begin
              _T_1259 <= _T_1265;
            end else begin
              _T_1259 <= _T_1256;
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1333 <= 1'h0;
    end else begin
      _T_1333 <= _T_1317;
    end
    if (_T_337) begin
      _T_1336 <= 2'h0;
    end else begin
      if (_T_1075) begin
        _T_1336 <= _T_1322;
      end
    end
    if (_T_337) begin
      _T_1339 <= 2'h0;
    end else begin
      if (_T_1075) begin
        _T_1339 <= _T_1007;
      end
    end
    if (_T_337) begin
      _T_1342 <= 1'h0;
    end else begin
      if (_T_1075) begin
        if (_T_1319) begin
          _T_1342 <= _T_1320;
        end else begin
          _T_1342 <= _T_985;
        end
      end
    end
    if (_T_337) begin
      _T_1345 <= 1'h0;
    end else begin
      if (_T_1075) begin
        _T_1345 <= _T_1108;
      end
    end
    if (_T_337) begin
      _T_1348 <= 1'h0;
    end else begin
      if (_T_1075) begin
        if (_T_959) begin
          _T_1348 <= 1'h1;
        end else begin
          if (_T_1072) begin
            _T_1348 <= 1'h0;
          end else begin
            _T_1348 <= _T_1052;
          end
        end
      end
    end
    if (_T_337) begin
      _T_1351 <= 2'h0;
    end else begin
      if (_T_1075) begin
        _T_1351 <= _T_984;
      end
    end
    if (_T_337) begin
      _T_1354 <= 1'h0;
    end else begin
      if (_T_1325) begin
        _T_1354 <= _T_959;
      end
    end
    if (_T_337) begin
      _T_1357 <= 9'h0;
    end else begin
      if (_T_1075) begin
        _T_1357 <= _T_1330;
      end
    end
    if (_T_337) begin
      _T_1360 <= 1'h0;
    end else begin
      if (_T_1075) begin
        _T_1360 <= _T_1362;
      end
    end
    if (_T_337) begin
      _T_1365 <= 13'h0;
    end else begin
      if (_T_1111) begin
        if (_T_347) begin
          _T_1365 <= 13'h0;
        end else begin
          if (_T_1390) begin
            _T_1365 <= 13'h0;
          end else begin
            _T_1365 <= _T_1393;
          end
        end
      end
    end
    if (_T_337) begin
      _T_1368 <= 13'h0;
    end else begin
      if (_T_1399) begin
        _T_1368 <= _T_1365;
      end
    end
    if (_T_337) begin
      _T_1371 <= 13'h0;
    end else begin
      if (_T_1432) begin
        _T_1371 <= _T_1401;
      end
    end
    if (_T_337) begin
      _T_1374 <= 13'h0;
    end else begin
      if (_T_1432) begin
        _T_1374 <= _T_1403;
      end
    end
    if (_T_337) begin
      _T_1377 <= 13'h0;
    end else begin
      if (_T_1432) begin
        _T_1377 <= _T_1405;
      end
    end
    if (_T_337) begin
      _T_1380 <= 13'h0;
    end else begin
      if (_T_1433) begin
        _T_1380 <= _T_1409;
      end
    end
    if (_T_337) begin
      _T_1383 <= 13'h0;
    end else begin
      _T_1383 <= _GEN_95[12:0];
    end
    if (_T_337) begin
      _T_1476_0 <= 13'h1fff;
    end else begin
      _T_1476_0 <= _GEN_96[12:0];
    end
    if (_T_337) begin
      _T_1476_1 <= 13'h1fff;
    end else begin
      _T_1476_1 <= _GEN_97[12:0];
    end
    if (_T_337) begin
      _T_1476_2 <= 13'h1fff;
    end else begin
      _T_1476_2 <= _GEN_98[12:0];
    end
    if (_T_337) begin
      _T_1476_3 <= 13'h1fff;
    end else begin
      _T_1476_3 <= _GEN_99[12:0];
    end
    if (_T_337) begin
      _T_1495 <= 1'h0;
    end else begin
      _T_1495 <= _T_1608;
    end
    if (_T_337) begin
      _T_1502 <= 15'h1fff;
    end else begin
      if (_T_1639) begin
        if (_T_1567) begin
          _T_1502 <= 15'h1fff;
        end else begin
          if (_T_1557) begin
            _T_1502 <= _T_1566;
          end else begin
            _T_1502 <= _T_1550;
          end
        end
      end
    end
    if (_T_337) begin
      _T_1505 <= 1'h0;
    end else begin
      _T_1505 <= _T_1049;
    end
    if (_T_337) begin
      _T_1511 <= 2'h0;
    end else begin
      if (_T_1052) begin
        _T_1511 <= _T_1336;
      end
    end
    if (_T_337) begin
      _T_1514 <= 2'h0;
    end else begin
      if (_T_1052) begin
        _T_1514 <= _T_1339;
      end
    end
    if (_T_337) begin
      _T_1517 <= 1'h0;
    end else begin
      if (_T_1052) begin
        _T_1517 <= _T_1342;
      end
    end
    if (_T_337) begin
      _T_1520 <= 1'h0;
    end else begin
      if (_T_1052) begin
        _T_1520 <= _T_1345;
      end
    end
    if (_T_337) begin
      _T_1523 <= 8'h0;
    end else begin
      if (_T_1052) begin
        _T_1523 <= _T_1078;
      end
    end
    if (_T_337) begin
      _T_1526 <= 1'h0;
    end else begin
      if (_T_1052) begin
        _T_1526 <= _T_1348;
      end
    end
    if (_T_337) begin
      _T_1529 <= 2'h0;
    end else begin
      if (_T_1052) begin
        _T_1529 <= _T_1351;
      end
    end
    if (_T_337) begin
      _T_1532 <= 1'h0;
    end else begin
      if (_T_1052) begin
        _T_1532 <= _T_1354;
      end
    end
    if (_T_337) begin
      _T_1535 <= 1'h0;
    end else begin
      if (_T_1052) begin
        _T_1535 <= _T_1360;
      end
    end
    if (_T_337) begin
      _T_1538 <= 9'h0;
    end else begin
      if (_T_1052) begin
        _T_1538 <= _T_1357;
      end else begin
        _T_1538 <= {{8'd0}, _T_1052};
      end
    end
    if (_T_337) begin
      _T_1660 <= 1'h0;
    end else begin
      _T_1660 <= _T_1505;
    end
    if (_T_337) begin
      _T_1663 <= 1'h0;
    end else begin
      _T_1663 <= _T_1660;
    end
    if (_T_337) begin
      _T_1666 <= 1'h0;
    end else begin
      _T_1666 <= _T_1663;
    end
    if (_T_337) begin
      _T_1669 <= 1'h0;
    end else begin
      _T_1669 <= _T_1666;
    end
    if (_T_337) begin
      _T_1672 <= 1'h0;
    end else begin
      _T_1672 <= _T_1669;
    end
    if (_T_337) begin
      _T_1675 <= 1'h0;
    end else begin
      _T_1675 <= _T_1672;
    end
    if (_T_337) begin
      _T_1680 <= 29'h0;
    end else begin
      if (_T_1505) begin
        _T_1680 <= _T_1655;
      end
    end
    if (_T_337) begin
      _T_1683 <= 29'h0;
    end else begin
      if (_T_1660) begin
        _T_1683 <= _T_1680;
      end
    end
    if (_T_337) begin
      _T_1686 <= 29'h0;
    end else begin
      if (_T_1663) begin
        _T_1686 <= _T_1683;
      end
    end
    if (_T_337) begin
      _T_1689 <= 29'h0;
    end else begin
      if (_T_1666) begin
        _T_1689 <= _T_1686;
      end
    end
    if (_T_337) begin
      _T_1692 <= 29'h0;
    end else begin
      if (_T_1669) begin
        _T_1692 <= _T_1689;
      end
    end
    if (_T_337) begin
      _T_1695 <= 29'h0;
    end else begin
      if (_T_1672) begin
        _T_1695 <= _T_1692;
      end
    end
    if (_T_337) begin
      _T_1768 <= 1'h1;
    end else begin
      if (sc2buf_dat_rd_valid) begin
        _T_1768 <= 1'h0;
      end
    end
    if (_T_337) begin
      _T_1780 <= 1'h1;
    end else begin
      if (_T_1825) begin
        _T_1780 <= 1'h0;
      end else begin
        if (sc2buf_dat_rd_valid) begin
          _T_1780 <= _T_1768;
        end
      end
    end
    if (sc2buf_dat_rd_valid) begin
      _T_1791 <= sc2buf_dat_rd_data;
    end
    if (_T_1825) begin
      _T_1799 <= _T_1791;
    end
    if (_T_337) begin
      _T_1899 <= 8'h0;
    end else begin
      if (_T_2105) begin
        if (_T_347) begin
          _T_1899 <= 8'h40;
        end else begin
          if (_T_2061) begin
            _T_1899 <= _T_1911;
          end else begin
            if (_T_2062) begin
              _T_1899 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1899 <= 8'h40;
              end else begin
                _T_1899 <= _T_2030;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1902 <= 8'h0;
    end else begin
      if (_T_2111) begin
        if (_T_347) begin
          _T_1902 <= 8'h40;
        end else begin
          if (_T_2072) begin
            _T_1902 <= _T_1914;
          end else begin
            if (_T_2073) begin
              _T_1902 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1902 <= 8'h40;
              end else begin
                _T_1902 <= _T_2039;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1905 <= 8'h0;
    end else begin
      if (_T_2117) begin
        if (_T_347) begin
          _T_1905 <= 8'h40;
        end else begin
          if (_T_2083) begin
            _T_1905 <= _T_1917;
          end else begin
            if (_T_2084) begin
              _T_1905 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1905 <= 8'h40;
              end else begin
                _T_1905 <= _T_2048;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1908 <= 8'h0;
    end else begin
      if (_T_2123) begin
        if (_T_347) begin
          _T_1908 <= 8'h40;
        end else begin
          if (_T_2094) begin
            _T_1908 <= _T_1920;
          end else begin
            if (_T_2095) begin
              _T_1908 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1908 <= 8'h40;
              end else begin
                _T_1908 <= _T_2057;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1911 <= 8'h0;
    end else begin
      if (_T_2128) begin
        if (_T_347) begin
          _T_1911 <= 8'h40;
        end else begin
          if (!(_T_2061)) begin
            if (_T_2062) begin
              _T_1911 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1911 <= 8'h40;
              end else begin
                _T_1911 <= _T_2030;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1914 <= 8'h0;
    end else begin
      if (_T_2136) begin
        if (_T_347) begin
          _T_1914 <= 8'h40;
        end else begin
          if (!(_T_2072)) begin
            if (_T_2073) begin
              _T_1914 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1914 <= 8'h40;
              end else begin
                _T_1914 <= _T_2039;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1917 <= 8'h0;
    end else begin
      if (_T_2144) begin
        if (_T_347) begin
          _T_1917 <= 8'h40;
        end else begin
          if (!(_T_2083)) begin
            if (_T_2084) begin
              _T_1917 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1917 <= 8'h40;
              end else begin
                _T_1917 <= _T_2048;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1920 <= 8'h0;
    end else begin
      if (_T_2152) begin
        if (_T_347) begin
          _T_1920 <= 8'h40;
        end else begin
          if (!(_T_2094)) begin
            if (_T_2095) begin
              _T_1920 <= 8'h40;
            end else begin
              if (_T_2024) begin
                _T_1920 <= 8'h40;
              end else begin
                _T_1920 <= _T_2057;
              end
            end
          end
        end
      end
    end
    if (_T_337) begin
      _T_1931 <= 1'h0;
    end else begin
      _T_1931 <= _T_1928;
    end
    if (_T_337) begin
      _T_1945 <= 27'h0;
    end else begin
      if (_T_1928) begin
        _T_1945 <= _T_1942;
      end
    end
    _T_2328 <= _GEN_149[255:0];
    _T_2330 <= _GEN_150[127:0];
    if (_T_2538) begin
      _T_2332 <= _T_2330;
    end
    _T_2334 <= _GEN_151[127:0];
    if (_T_2538) begin
      _T_2336 <= _T_2334;
    end
    _T_2338 <= _GEN_154[127:0];
    if (_T_337) begin
      _T_3136 <= 1'h0;
    end else begin
      _T_3136 <= _T_1965;
    end
    if (_T_337) begin
      _T_3406_0 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_0 <= _T_2937;
      end
    end
    if (_T_337) begin
      _T_3406_1 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_1 <= _T_2939;
      end
    end
    if (_T_337) begin
      _T_3406_2 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_2 <= _T_2941;
      end
    end
    if (_T_337) begin
      _T_3406_3 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_3 <= _T_2943;
      end
    end
    if (_T_337) begin
      _T_3406_4 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_4 <= _T_2945;
      end
    end
    if (_T_337) begin
      _T_3406_5 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_5 <= _T_2947;
      end
    end
    if (_T_337) begin
      _T_3406_6 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_6 <= _T_2949;
      end
    end
    if (_T_337) begin
      _T_3406_7 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_7 <= _T_2951;
      end
    end
    if (_T_337) begin
      _T_3406_8 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_8 <= _T_2953;
      end
    end
    if (_T_337) begin
      _T_3406_9 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_9 <= _T_2955;
      end
    end
    if (_T_337) begin
      _T_3406_10 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_10 <= _T_2957;
      end
    end
    if (_T_337) begin
      _T_3406_11 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_11 <= _T_2959;
      end
    end
    if (_T_337) begin
      _T_3406_12 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_12 <= _T_2961;
      end
    end
    if (_T_337) begin
      _T_3406_13 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_13 <= _T_2963;
      end
    end
    if (_T_337) begin
      _T_3406_14 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_14 <= _T_2965;
      end
    end
    if (_T_337) begin
      _T_3406_15 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_15 <= _T_2967;
      end
    end
    if (_T_337) begin
      _T_3406_16 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_16 <= _T_2969;
      end
    end
    if (_T_337) begin
      _T_3406_17 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_17 <= _T_2971;
      end
    end
    if (_T_337) begin
      _T_3406_18 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_18 <= _T_2973;
      end
    end
    if (_T_337) begin
      _T_3406_19 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_19 <= _T_2975;
      end
    end
    if (_T_337) begin
      _T_3406_20 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_20 <= _T_2977;
      end
    end
    if (_T_337) begin
      _T_3406_21 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_21 <= _T_2979;
      end
    end
    if (_T_337) begin
      _T_3406_22 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_22 <= _T_2981;
      end
    end
    if (_T_337) begin
      _T_3406_23 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_23 <= _T_2983;
      end
    end
    if (_T_337) begin
      _T_3406_24 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_24 <= _T_2985;
      end
    end
    if (_T_337) begin
      _T_3406_25 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_25 <= _T_2987;
      end
    end
    if (_T_337) begin
      _T_3406_26 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_26 <= _T_2989;
      end
    end
    if (_T_337) begin
      _T_3406_27 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_27 <= _T_2991;
      end
    end
    if (_T_337) begin
      _T_3406_28 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_28 <= _T_2993;
      end
    end
    if (_T_337) begin
      _T_3406_29 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_29 <= _T_2995;
      end
    end
    if (_T_337) begin
      _T_3406_30 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_30 <= _T_2997;
      end
    end
    if (_T_337) begin
      _T_3406_31 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_31 <= _T_2999;
      end
    end
    if (_T_337) begin
      _T_3406_32 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_32 <= _T_3001;
      end
    end
    if (_T_337) begin
      _T_3406_33 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_33 <= _T_3003;
      end
    end
    if (_T_337) begin
      _T_3406_34 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_34 <= _T_3005;
      end
    end
    if (_T_337) begin
      _T_3406_35 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_35 <= _T_3007;
      end
    end
    if (_T_337) begin
      _T_3406_36 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_36 <= _T_3009;
      end
    end
    if (_T_337) begin
      _T_3406_37 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_37 <= _T_3011;
      end
    end
    if (_T_337) begin
      _T_3406_38 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_38 <= _T_3013;
      end
    end
    if (_T_337) begin
      _T_3406_39 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_39 <= _T_3015;
      end
    end
    if (_T_337) begin
      _T_3406_40 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_40 <= _T_3017;
      end
    end
    if (_T_337) begin
      _T_3406_41 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_41 <= _T_3019;
      end
    end
    if (_T_337) begin
      _T_3406_42 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_42 <= _T_3021;
      end
    end
    if (_T_337) begin
      _T_3406_43 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_43 <= _T_3023;
      end
    end
    if (_T_337) begin
      _T_3406_44 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_44 <= _T_3025;
      end
    end
    if (_T_337) begin
      _T_3406_45 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_45 <= _T_3027;
      end
    end
    if (_T_337) begin
      _T_3406_46 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_46 <= _T_3029;
      end
    end
    if (_T_337) begin
      _T_3406_47 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_47 <= _T_3031;
      end
    end
    if (_T_337) begin
      _T_3406_48 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_48 <= _T_3033;
      end
    end
    if (_T_337) begin
      _T_3406_49 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_49 <= _T_3035;
      end
    end
    if (_T_337) begin
      _T_3406_50 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_50 <= _T_3037;
      end
    end
    if (_T_337) begin
      _T_3406_51 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_51 <= _T_3039;
      end
    end
    if (_T_337) begin
      _T_3406_52 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_52 <= _T_3041;
      end
    end
    if (_T_337) begin
      _T_3406_53 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_53 <= _T_3043;
      end
    end
    if (_T_337) begin
      _T_3406_54 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_54 <= _T_3045;
      end
    end
    if (_T_337) begin
      _T_3406_55 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_55 <= _T_3047;
      end
    end
    if (_T_337) begin
      _T_3406_56 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_56 <= _T_3049;
      end
    end
    if (_T_337) begin
      _T_3406_57 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_57 <= _T_3051;
      end
    end
    if (_T_337) begin
      _T_3406_58 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_58 <= _T_3053;
      end
    end
    if (_T_337) begin
      _T_3406_59 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_59 <= _T_3055;
      end
    end
    if (_T_337) begin
      _T_3406_60 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_60 <= _T_3057;
      end
    end
    if (_T_337) begin
      _T_3406_61 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_61 <= _T_3059;
      end
    end
    if (_T_337) begin
      _T_3406_62 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_62 <= _T_3061;
      end
    end
    if (_T_337) begin
      _T_3406_63 <= 1'h0;
    end else begin
      if (_T_1965) begin
        _T_3406_63 <= _T_3063;
      end
    end
    if (_T_3673) begin
      if (_T_2605) begin
        _T_3606_0 <= _T_2466;
      end else begin
        _T_3606_0 <= _T_2263;
      end
    end
    if (_T_3674) begin
      if (_T_2605) begin
        _T_3606_1 <= _T_2467;
      end else begin
        _T_3606_1 <= _T_2264;
      end
    end
    if (_T_3675) begin
      if (_T_2605) begin
        _T_3606_2 <= _T_2468;
      end else begin
        _T_3606_2 <= _T_2265;
      end
    end
    if (_T_3676) begin
      if (_T_2605) begin
        _T_3606_3 <= _T_2469;
      end else begin
        _T_3606_3 <= _T_2266;
      end
    end
    if (_T_3677) begin
      if (_T_2605) begin
        _T_3606_4 <= _T_2470;
      end else begin
        _T_3606_4 <= _T_2267;
      end
    end
    if (_T_3678) begin
      if (_T_2605) begin
        _T_3606_5 <= _T_2471;
      end else begin
        _T_3606_5 <= _T_2268;
      end
    end
    if (_T_3679) begin
      if (_T_2605) begin
        _T_3606_6 <= _T_2472;
      end else begin
        _T_3606_6 <= _T_2269;
      end
    end
    if (_T_3680) begin
      if (_T_2605) begin
        _T_3606_7 <= _T_2473;
      end else begin
        _T_3606_7 <= _T_2270;
      end
    end
    if (_T_3681) begin
      if (_T_2605) begin
        _T_3606_8 <= _T_2474;
      end else begin
        _T_3606_8 <= _T_2271;
      end
    end
    if (_T_3682) begin
      if (_T_2605) begin
        _T_3606_9 <= _T_2475;
      end else begin
        _T_3606_9 <= _T_2272;
      end
    end
    if (_T_3683) begin
      if (_T_2605) begin
        _T_3606_10 <= _T_2476;
      end else begin
        _T_3606_10 <= _T_2273;
      end
    end
    if (_T_3684) begin
      if (_T_2605) begin
        _T_3606_11 <= _T_2477;
      end else begin
        _T_3606_11 <= _T_2274;
      end
    end
    if (_T_3685) begin
      if (_T_2605) begin
        _T_3606_12 <= _T_2478;
      end else begin
        _T_3606_12 <= _T_2275;
      end
    end
    if (_T_3686) begin
      if (_T_2605) begin
        _T_3606_13 <= _T_2479;
      end else begin
        _T_3606_13 <= _T_2276;
      end
    end
    if (_T_3687) begin
      if (_T_2605) begin
        _T_3606_14 <= _T_2480;
      end else begin
        _T_3606_14 <= _T_2277;
      end
    end
    if (_T_3688) begin
      if (_T_2605) begin
        _T_3606_15 <= _T_2481;
      end else begin
        _T_3606_15 <= _T_2278;
      end
    end
    if (_T_3689) begin
      if (_T_2605) begin
        _T_3606_16 <= _T_2482;
      end else begin
        _T_3606_16 <= _T_2279;
      end
    end
    if (_T_3690) begin
      if (_T_2605) begin
        _T_3606_17 <= _T_2483;
      end else begin
        _T_3606_17 <= _T_2280;
      end
    end
    if (_T_3691) begin
      if (_T_2605) begin
        _T_3606_18 <= _T_2484;
      end else begin
        _T_3606_18 <= _T_2281;
      end
    end
    if (_T_3692) begin
      if (_T_2605) begin
        _T_3606_19 <= _T_2485;
      end else begin
        _T_3606_19 <= _T_2282;
      end
    end
    if (_T_3693) begin
      if (_T_2605) begin
        _T_3606_20 <= _T_2486;
      end else begin
        _T_3606_20 <= _T_2283;
      end
    end
    if (_T_3694) begin
      if (_T_2605) begin
        _T_3606_21 <= _T_2487;
      end else begin
        _T_3606_21 <= _T_2284;
      end
    end
    if (_T_3695) begin
      if (_T_2605) begin
        _T_3606_22 <= _T_2488;
      end else begin
        _T_3606_22 <= _T_2285;
      end
    end
    if (_T_3696) begin
      if (_T_2605) begin
        _T_3606_23 <= _T_2489;
      end else begin
        _T_3606_23 <= _T_2286;
      end
    end
    if (_T_3697) begin
      if (_T_2605) begin
        _T_3606_24 <= _T_2490;
      end else begin
        _T_3606_24 <= _T_2287;
      end
    end
    if (_T_3698) begin
      if (_T_2605) begin
        _T_3606_25 <= _T_2491;
      end else begin
        _T_3606_25 <= _T_2288;
      end
    end
    if (_T_3699) begin
      if (_T_2605) begin
        _T_3606_26 <= _T_2492;
      end else begin
        _T_3606_26 <= _T_2289;
      end
    end
    if (_T_3700) begin
      if (_T_2605) begin
        _T_3606_27 <= _T_2493;
      end else begin
        _T_3606_27 <= _T_2290;
      end
    end
    if (_T_3701) begin
      if (_T_2605) begin
        _T_3606_28 <= _T_2494;
      end else begin
        _T_3606_28 <= _T_2291;
      end
    end
    if (_T_3702) begin
      if (_T_2605) begin
        _T_3606_29 <= _T_2495;
      end else begin
        _T_3606_29 <= _T_2292;
      end
    end
    if (_T_3703) begin
      if (_T_2605) begin
        _T_3606_30 <= _T_2496;
      end else begin
        _T_3606_30 <= _T_2293;
      end
    end
    if (_T_3704) begin
      if (_T_2605) begin
        _T_3606_31 <= _T_2497;
      end else begin
        _T_3606_31 <= _T_2294;
      end
    end
    if (_T_3705) begin
      if (_T_2605) begin
        _T_3606_32 <= _T_2498;
      end else begin
        _T_3606_32 <= _T_2295;
      end
    end
    if (_T_3706) begin
      if (_T_2605) begin
        _T_3606_33 <= _T_2499;
      end else begin
        _T_3606_33 <= _T_2296;
      end
    end
    if (_T_3707) begin
      if (_T_2605) begin
        _T_3606_34 <= _T_2500;
      end else begin
        _T_3606_34 <= _T_2297;
      end
    end
    if (_T_3708) begin
      if (_T_2605) begin
        _T_3606_35 <= _T_2501;
      end else begin
        _T_3606_35 <= _T_2298;
      end
    end
    if (_T_3709) begin
      if (_T_2605) begin
        _T_3606_36 <= _T_2502;
      end else begin
        _T_3606_36 <= _T_2299;
      end
    end
    if (_T_3710) begin
      if (_T_2605) begin
        _T_3606_37 <= _T_2503;
      end else begin
        _T_3606_37 <= _T_2300;
      end
    end
    if (_T_3711) begin
      if (_T_2605) begin
        _T_3606_38 <= _T_2504;
      end else begin
        _T_3606_38 <= _T_2301;
      end
    end
    if (_T_3712) begin
      if (_T_2605) begin
        _T_3606_39 <= _T_2505;
      end else begin
        _T_3606_39 <= _T_2302;
      end
    end
    if (_T_3713) begin
      if (_T_2605) begin
        _T_3606_40 <= _T_2506;
      end else begin
        _T_3606_40 <= _T_2303;
      end
    end
    if (_T_3714) begin
      if (_T_2605) begin
        _T_3606_41 <= _T_2507;
      end else begin
        _T_3606_41 <= _T_2304;
      end
    end
    if (_T_3715) begin
      if (_T_2605) begin
        _T_3606_42 <= _T_2508;
      end else begin
        _T_3606_42 <= _T_2305;
      end
    end
    if (_T_3716) begin
      if (_T_2605) begin
        _T_3606_43 <= _T_2509;
      end else begin
        _T_3606_43 <= _T_2306;
      end
    end
    if (_T_3717) begin
      if (_T_2605) begin
        _T_3606_44 <= _T_2510;
      end else begin
        _T_3606_44 <= _T_2307;
      end
    end
    if (_T_3718) begin
      if (_T_2605) begin
        _T_3606_45 <= _T_2511;
      end else begin
        _T_3606_45 <= _T_2308;
      end
    end
    if (_T_3719) begin
      if (_T_2605) begin
        _T_3606_46 <= _T_2512;
      end else begin
        _T_3606_46 <= _T_2309;
      end
    end
    if (_T_3720) begin
      if (_T_2605) begin
        _T_3606_47 <= _T_2513;
      end else begin
        _T_3606_47 <= _T_2310;
      end
    end
    if (_T_3721) begin
      if (_T_2605) begin
        _T_3606_48 <= _T_2514;
      end else begin
        _T_3606_48 <= _T_2311;
      end
    end
    if (_T_3722) begin
      if (_T_2605) begin
        _T_3606_49 <= _T_2515;
      end else begin
        _T_3606_49 <= _T_2312;
      end
    end
    if (_T_3723) begin
      if (_T_2605) begin
        _T_3606_50 <= _T_2516;
      end else begin
        _T_3606_50 <= _T_2313;
      end
    end
    if (_T_3724) begin
      if (_T_2605) begin
        _T_3606_51 <= _T_2517;
      end else begin
        _T_3606_51 <= _T_2314;
      end
    end
    if (_T_3725) begin
      if (_T_2605) begin
        _T_3606_52 <= _T_2518;
      end else begin
        _T_3606_52 <= _T_2315;
      end
    end
    if (_T_3726) begin
      if (_T_2605) begin
        _T_3606_53 <= _T_2519;
      end else begin
        _T_3606_53 <= _T_2316;
      end
    end
    if (_T_3727) begin
      if (_T_2605) begin
        _T_3606_54 <= _T_2520;
      end else begin
        _T_3606_54 <= _T_2317;
      end
    end
    if (_T_3728) begin
      if (_T_2605) begin
        _T_3606_55 <= _T_2521;
      end else begin
        _T_3606_55 <= _T_2318;
      end
    end
    if (_T_3729) begin
      if (_T_2605) begin
        _T_3606_56 <= _T_2522;
      end else begin
        _T_3606_56 <= _T_2319;
      end
    end
    if (_T_3730) begin
      if (_T_2605) begin
        _T_3606_57 <= _T_2523;
      end else begin
        _T_3606_57 <= _T_2320;
      end
    end
    if (_T_3731) begin
      if (_T_2605) begin
        _T_3606_58 <= _T_2524;
      end else begin
        _T_3606_58 <= _T_2321;
      end
    end
    if (_T_3732) begin
      if (_T_2605) begin
        _T_3606_59 <= _T_2525;
      end else begin
        _T_3606_59 <= _T_2322;
      end
    end
    if (_T_3733) begin
      if (_T_2605) begin
        _T_3606_60 <= _T_2526;
      end else begin
        _T_3606_60 <= _T_2323;
      end
    end
    if (_T_3734) begin
      if (_T_2605) begin
        _T_3606_61 <= _T_2527;
      end else begin
        _T_3606_61 <= _T_2324;
      end
    end
    if (_T_3735) begin
      if (_T_2605) begin
        _T_3606_62 <= _T_2528;
      end else begin
        _T_3606_62 <= _T_2325;
      end
    end
    if (_T_3736) begin
      if (_T_2605) begin
        _T_3606_63 <= _T_2529;
      end else begin
        _T_3606_63 <= _T_2326;
      end
    end
    if (_T_337) begin
      _T_3739 <= 1'h0;
    end else begin
      _T_3739 <= _T_3136;
    end
    if (_T_337) begin
      _T_4006_0 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_0 <= 1'h0;
        end else begin
          _T_4006_0 <= _T_3406_0;
        end
      end
    end
    if (_T_337) begin
      _T_4006_1 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_1 <= 1'h0;
        end else begin
          _T_4006_1 <= _T_3406_1;
        end
      end
    end
    if (_T_337) begin
      _T_4006_2 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_2 <= 1'h0;
        end else begin
          _T_4006_2 <= _T_3406_2;
        end
      end
    end
    if (_T_337) begin
      _T_4006_3 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_3 <= 1'h0;
        end else begin
          _T_4006_3 <= _T_3406_3;
        end
      end
    end
    if (_T_337) begin
      _T_4006_4 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_4 <= 1'h0;
        end else begin
          _T_4006_4 <= _T_3406_4;
        end
      end
    end
    if (_T_337) begin
      _T_4006_5 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_5 <= 1'h0;
        end else begin
          _T_4006_5 <= _T_3406_5;
        end
      end
    end
    if (_T_337) begin
      _T_4006_6 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_6 <= 1'h0;
        end else begin
          _T_4006_6 <= _T_3406_6;
        end
      end
    end
    if (_T_337) begin
      _T_4006_7 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_7 <= 1'h0;
        end else begin
          _T_4006_7 <= _T_3406_7;
        end
      end
    end
    if (_T_337) begin
      _T_4006_8 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_8 <= 1'h0;
        end else begin
          _T_4006_8 <= _T_3406_8;
        end
      end
    end
    if (_T_337) begin
      _T_4006_9 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_9 <= 1'h0;
        end else begin
          _T_4006_9 <= _T_3406_9;
        end
      end
    end
    if (_T_337) begin
      _T_4006_10 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_10 <= 1'h0;
        end else begin
          _T_4006_10 <= _T_3406_10;
        end
      end
    end
    if (_T_337) begin
      _T_4006_11 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_11 <= 1'h0;
        end else begin
          _T_4006_11 <= _T_3406_11;
        end
      end
    end
    if (_T_337) begin
      _T_4006_12 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_12 <= 1'h0;
        end else begin
          _T_4006_12 <= _T_3406_12;
        end
      end
    end
    if (_T_337) begin
      _T_4006_13 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_13 <= 1'h0;
        end else begin
          _T_4006_13 <= _T_3406_13;
        end
      end
    end
    if (_T_337) begin
      _T_4006_14 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_14 <= 1'h0;
        end else begin
          _T_4006_14 <= _T_3406_14;
        end
      end
    end
    if (_T_337) begin
      _T_4006_15 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_15 <= 1'h0;
        end else begin
          _T_4006_15 <= _T_3406_15;
        end
      end
    end
    if (_T_337) begin
      _T_4006_16 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_16 <= 1'h0;
        end else begin
          _T_4006_16 <= _T_3406_16;
        end
      end
    end
    if (_T_337) begin
      _T_4006_17 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_17 <= 1'h0;
        end else begin
          _T_4006_17 <= _T_3406_17;
        end
      end
    end
    if (_T_337) begin
      _T_4006_18 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_18 <= 1'h0;
        end else begin
          _T_4006_18 <= _T_3406_18;
        end
      end
    end
    if (_T_337) begin
      _T_4006_19 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_19 <= 1'h0;
        end else begin
          _T_4006_19 <= _T_3406_19;
        end
      end
    end
    if (_T_337) begin
      _T_4006_20 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_20 <= 1'h0;
        end else begin
          _T_4006_20 <= _T_3406_20;
        end
      end
    end
    if (_T_337) begin
      _T_4006_21 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_21 <= 1'h0;
        end else begin
          _T_4006_21 <= _T_3406_21;
        end
      end
    end
    if (_T_337) begin
      _T_4006_22 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_22 <= 1'h0;
        end else begin
          _T_4006_22 <= _T_3406_22;
        end
      end
    end
    if (_T_337) begin
      _T_4006_23 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_23 <= 1'h0;
        end else begin
          _T_4006_23 <= _T_3406_23;
        end
      end
    end
    if (_T_337) begin
      _T_4006_24 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_24 <= 1'h0;
        end else begin
          _T_4006_24 <= _T_3406_24;
        end
      end
    end
    if (_T_337) begin
      _T_4006_25 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_25 <= 1'h0;
        end else begin
          _T_4006_25 <= _T_3406_25;
        end
      end
    end
    if (_T_337) begin
      _T_4006_26 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_26 <= 1'h0;
        end else begin
          _T_4006_26 <= _T_3406_26;
        end
      end
    end
    if (_T_337) begin
      _T_4006_27 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_27 <= 1'h0;
        end else begin
          _T_4006_27 <= _T_3406_27;
        end
      end
    end
    if (_T_337) begin
      _T_4006_28 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_28 <= 1'h0;
        end else begin
          _T_4006_28 <= _T_3406_28;
        end
      end
    end
    if (_T_337) begin
      _T_4006_29 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_29 <= 1'h0;
        end else begin
          _T_4006_29 <= _T_3406_29;
        end
      end
    end
    if (_T_337) begin
      _T_4006_30 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_30 <= 1'h0;
        end else begin
          _T_4006_30 <= _T_3406_30;
        end
      end
    end
    if (_T_337) begin
      _T_4006_31 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_31 <= 1'h0;
        end else begin
          _T_4006_31 <= _T_3406_31;
        end
      end
    end
    if (_T_337) begin
      _T_4006_32 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_32 <= 1'h0;
        end else begin
          _T_4006_32 <= _T_3406_32;
        end
      end
    end
    if (_T_337) begin
      _T_4006_33 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_33 <= 1'h0;
        end else begin
          _T_4006_33 <= _T_3406_33;
        end
      end
    end
    if (_T_337) begin
      _T_4006_34 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_34 <= 1'h0;
        end else begin
          _T_4006_34 <= _T_3406_34;
        end
      end
    end
    if (_T_337) begin
      _T_4006_35 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_35 <= 1'h0;
        end else begin
          _T_4006_35 <= _T_3406_35;
        end
      end
    end
    if (_T_337) begin
      _T_4006_36 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_36 <= 1'h0;
        end else begin
          _T_4006_36 <= _T_3406_36;
        end
      end
    end
    if (_T_337) begin
      _T_4006_37 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_37 <= 1'h0;
        end else begin
          _T_4006_37 <= _T_3406_37;
        end
      end
    end
    if (_T_337) begin
      _T_4006_38 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_38 <= 1'h0;
        end else begin
          _T_4006_38 <= _T_3406_38;
        end
      end
    end
    if (_T_337) begin
      _T_4006_39 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_39 <= 1'h0;
        end else begin
          _T_4006_39 <= _T_3406_39;
        end
      end
    end
    if (_T_337) begin
      _T_4006_40 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_40 <= 1'h0;
        end else begin
          _T_4006_40 <= _T_3406_40;
        end
      end
    end
    if (_T_337) begin
      _T_4006_41 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_41 <= 1'h0;
        end else begin
          _T_4006_41 <= _T_3406_41;
        end
      end
    end
    if (_T_337) begin
      _T_4006_42 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_42 <= 1'h0;
        end else begin
          _T_4006_42 <= _T_3406_42;
        end
      end
    end
    if (_T_337) begin
      _T_4006_43 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_43 <= 1'h0;
        end else begin
          _T_4006_43 <= _T_3406_43;
        end
      end
    end
    if (_T_337) begin
      _T_4006_44 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_44 <= 1'h0;
        end else begin
          _T_4006_44 <= _T_3406_44;
        end
      end
    end
    if (_T_337) begin
      _T_4006_45 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_45 <= 1'h0;
        end else begin
          _T_4006_45 <= _T_3406_45;
        end
      end
    end
    if (_T_337) begin
      _T_4006_46 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_46 <= 1'h0;
        end else begin
          _T_4006_46 <= _T_3406_46;
        end
      end
    end
    if (_T_337) begin
      _T_4006_47 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_47 <= 1'h0;
        end else begin
          _T_4006_47 <= _T_3406_47;
        end
      end
    end
    if (_T_337) begin
      _T_4006_48 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_48 <= 1'h0;
        end else begin
          _T_4006_48 <= _T_3406_48;
        end
      end
    end
    if (_T_337) begin
      _T_4006_49 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_49 <= 1'h0;
        end else begin
          _T_4006_49 <= _T_3406_49;
        end
      end
    end
    if (_T_337) begin
      _T_4006_50 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_50 <= 1'h0;
        end else begin
          _T_4006_50 <= _T_3406_50;
        end
      end
    end
    if (_T_337) begin
      _T_4006_51 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_51 <= 1'h0;
        end else begin
          _T_4006_51 <= _T_3406_51;
        end
      end
    end
    if (_T_337) begin
      _T_4006_52 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_52 <= 1'h0;
        end else begin
          _T_4006_52 <= _T_3406_52;
        end
      end
    end
    if (_T_337) begin
      _T_4006_53 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_53 <= 1'h0;
        end else begin
          _T_4006_53 <= _T_3406_53;
        end
      end
    end
    if (_T_337) begin
      _T_4006_54 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_54 <= 1'h0;
        end else begin
          _T_4006_54 <= _T_3406_54;
        end
      end
    end
    if (_T_337) begin
      _T_4006_55 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_55 <= 1'h0;
        end else begin
          _T_4006_55 <= _T_3406_55;
        end
      end
    end
    if (_T_337) begin
      _T_4006_56 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_56 <= 1'h0;
        end else begin
          _T_4006_56 <= _T_3406_56;
        end
      end
    end
    if (_T_337) begin
      _T_4006_57 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_57 <= 1'h0;
        end else begin
          _T_4006_57 <= _T_3406_57;
        end
      end
    end
    if (_T_337) begin
      _T_4006_58 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_58 <= 1'h0;
        end else begin
          _T_4006_58 <= _T_3406_58;
        end
      end
    end
    if (_T_337) begin
      _T_4006_59 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_59 <= 1'h0;
        end else begin
          _T_4006_59 <= _T_3406_59;
        end
      end
    end
    if (_T_337) begin
      _T_4006_60 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_60 <= 1'h0;
        end else begin
          _T_4006_60 <= _T_3406_60;
        end
      end
    end
    if (_T_337) begin
      _T_4006_61 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_61 <= 1'h0;
        end else begin
          _T_4006_61 <= _T_3406_61;
        end
      end
    end
    if (_T_337) begin
      _T_4006_62 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_62 <= 1'h0;
        end else begin
          _T_4006_62 <= _T_3406_62;
        end
      end
    end
    if (_T_337) begin
      _T_4006_63 <= 1'h0;
    end else begin
      if (_T_4543) begin
        if (_T_4276) begin
          _T_4006_63 <= 1'h0;
        end else begin
          _T_4006_63 <= _T_3406_63;
        end
      end
    end
    if (_T_337) begin
      _T_4205 <= 9'h0;
    end else begin
      if (_T_3136) begin
        _T_4205 <= {{8'd0}, _T_3136};
      end
    end
    if (_T_4411_0) begin
      _T_4209_0 <= _T_3606_0;
    end
    if (_T_4411_1) begin
      _T_4209_1 <= _T_3606_1;
    end
    if (_T_4411_2) begin
      _T_4209_2 <= _T_3606_2;
    end
    if (_T_4411_3) begin
      _T_4209_3 <= _T_3606_3;
    end
    if (_T_4411_4) begin
      _T_4209_4 <= _T_3606_4;
    end
    if (_T_4411_5) begin
      _T_4209_5 <= _T_3606_5;
    end
    if (_T_4411_6) begin
      _T_4209_6 <= _T_3606_6;
    end
    if (_T_4411_7) begin
      _T_4209_7 <= _T_3606_7;
    end
    if (_T_4411_8) begin
      _T_4209_8 <= _T_3606_8;
    end
    if (_T_4411_9) begin
      _T_4209_9 <= _T_3606_9;
    end
    if (_T_4411_10) begin
      _T_4209_10 <= _T_3606_10;
    end
    if (_T_4411_11) begin
      _T_4209_11 <= _T_3606_11;
    end
    if (_T_4411_12) begin
      _T_4209_12 <= _T_3606_12;
    end
    if (_T_4411_13) begin
      _T_4209_13 <= _T_3606_13;
    end
    if (_T_4411_14) begin
      _T_4209_14 <= _T_3606_14;
    end
    if (_T_4411_15) begin
      _T_4209_15 <= _T_3606_15;
    end
    if (_T_4411_16) begin
      _T_4209_16 <= _T_3606_16;
    end
    if (_T_4411_17) begin
      _T_4209_17 <= _T_3606_17;
    end
    if (_T_4411_18) begin
      _T_4209_18 <= _T_3606_18;
    end
    if (_T_4411_19) begin
      _T_4209_19 <= _T_3606_19;
    end
    if (_T_4411_20) begin
      _T_4209_20 <= _T_3606_20;
    end
    if (_T_4411_21) begin
      _T_4209_21 <= _T_3606_21;
    end
    if (_T_4411_22) begin
      _T_4209_22 <= _T_3606_22;
    end
    if (_T_4411_23) begin
      _T_4209_23 <= _T_3606_23;
    end
    if (_T_4411_24) begin
      _T_4209_24 <= _T_3606_24;
    end
    if (_T_4411_25) begin
      _T_4209_25 <= _T_3606_25;
    end
    if (_T_4411_26) begin
      _T_4209_26 <= _T_3606_26;
    end
    if (_T_4411_27) begin
      _T_4209_27 <= _T_3606_27;
    end
    if (_T_4411_28) begin
      _T_4209_28 <= _T_3606_28;
    end
    if (_T_4411_29) begin
      _T_4209_29 <= _T_3606_29;
    end
    if (_T_4411_30) begin
      _T_4209_30 <= _T_3606_30;
    end
    if (_T_4411_31) begin
      _T_4209_31 <= _T_3606_31;
    end
    if (_T_4411_32) begin
      _T_4209_32 <= _T_3606_32;
    end
    if (_T_4411_33) begin
      _T_4209_33 <= _T_3606_33;
    end
    if (_T_4411_34) begin
      _T_4209_34 <= _T_3606_34;
    end
    if (_T_4411_35) begin
      _T_4209_35 <= _T_3606_35;
    end
    if (_T_4411_36) begin
      _T_4209_36 <= _T_3606_36;
    end
    if (_T_4411_37) begin
      _T_4209_37 <= _T_3606_37;
    end
    if (_T_4411_38) begin
      _T_4209_38 <= _T_3606_38;
    end
    if (_T_4411_39) begin
      _T_4209_39 <= _T_3606_39;
    end
    if (_T_4411_40) begin
      _T_4209_40 <= _T_3606_40;
    end
    if (_T_4411_41) begin
      _T_4209_41 <= _T_3606_41;
    end
    if (_T_4411_42) begin
      _T_4209_42 <= _T_3606_42;
    end
    if (_T_4411_43) begin
      _T_4209_43 <= _T_3606_43;
    end
    if (_T_4411_44) begin
      _T_4209_44 <= _T_3606_44;
    end
    if (_T_4411_45) begin
      _T_4209_45 <= _T_3606_45;
    end
    if (_T_4411_46) begin
      _T_4209_46 <= _T_3606_46;
    end
    if (_T_4411_47) begin
      _T_4209_47 <= _T_3606_47;
    end
    if (_T_4411_48) begin
      _T_4209_48 <= _T_3606_48;
    end
    if (_T_4411_49) begin
      _T_4209_49 <= _T_3606_49;
    end
    if (_T_4411_50) begin
      _T_4209_50 <= _T_3606_50;
    end
    if (_T_4411_51) begin
      _T_4209_51 <= _T_3606_51;
    end
    if (_T_4411_52) begin
      _T_4209_52 <= _T_3606_52;
    end
    if (_T_4411_53) begin
      _T_4209_53 <= _T_3606_53;
    end
    if (_T_4411_54) begin
      _T_4209_54 <= _T_3606_54;
    end
    if (_T_4411_55) begin
      _T_4209_55 <= _T_3606_55;
    end
    if (_T_4411_56) begin
      _T_4209_56 <= _T_3606_56;
    end
    if (_T_4411_57) begin
      _T_4209_57 <= _T_3606_57;
    end
    if (_T_4411_58) begin
      _T_4209_58 <= _T_3606_58;
    end
    if (_T_4411_59) begin
      _T_4209_59 <= _T_3606_59;
    end
    if (_T_4411_60) begin
      _T_4209_60 <= _T_3606_60;
    end
    if (_T_4411_61) begin
      _T_4209_61 <= _T_3606_61;
    end
    if (_T_4411_62) begin
      _T_4209_62 <= _T_3606_62;
    end
    if (_T_4411_63) begin
      _T_4209_63 <= _T_3606_63;
    end
    if (_T_337) begin
      _T_4546 <= 1'h0;
    end else begin
      _T_4546 <= _T_3739;
    end
    if (_T_337) begin
      _T_4552 <= 1'h0;
    end else begin
      _T_4552 <= _T_3739;
    end
    if (_T_337) begin
      _T_4555 <= 1'h0;
    end else begin
      _T_4555 <= _T_3739;
    end
    if (_T_337) begin
      _T_4559 <= 9'h0;
    end else begin
      if (_T_4557) begin
        if (_T_4547) begin
          _T_4559 <= 9'h0;
        end else begin
          _T_4559 <= _T_4205;
        end
      end
    end
    if (_T_337) begin
      _T_4563 <= 9'h0;
    end else begin
      if (_T_4557) begin
        if (_T_4547) begin
          _T_4563 <= 9'h0;
        end else begin
          _T_4563 <= _T_4205;
        end
      end
    end
    if (_T_337) begin
      _T_4831_0 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_0 <= _T_4006_0;
      end
    end
    if (_T_337) begin
      _T_4831_1 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_1 <= _T_4006_1;
      end
    end
    if (_T_337) begin
      _T_4831_2 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_2 <= _T_4006_2;
      end
    end
    if (_T_337) begin
      _T_4831_3 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_3 <= _T_4006_3;
      end
    end
    if (_T_337) begin
      _T_4831_4 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_4 <= _T_4006_4;
      end
    end
    if (_T_337) begin
      _T_4831_5 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_5 <= _T_4006_5;
      end
    end
    if (_T_337) begin
      _T_4831_6 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_6 <= _T_4006_6;
      end
    end
    if (_T_337) begin
      _T_4831_7 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_7 <= _T_4006_7;
      end
    end
    if (_T_337) begin
      _T_4831_8 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_8 <= _T_4006_8;
      end
    end
    if (_T_337) begin
      _T_4831_9 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_9 <= _T_4006_9;
      end
    end
    if (_T_337) begin
      _T_4831_10 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_10 <= _T_4006_10;
      end
    end
    if (_T_337) begin
      _T_4831_11 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_11 <= _T_4006_11;
      end
    end
    if (_T_337) begin
      _T_4831_12 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_12 <= _T_4006_12;
      end
    end
    if (_T_337) begin
      _T_4831_13 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_13 <= _T_4006_13;
      end
    end
    if (_T_337) begin
      _T_4831_14 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_14 <= _T_4006_14;
      end
    end
    if (_T_337) begin
      _T_4831_15 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_15 <= _T_4006_15;
      end
    end
    if (_T_337) begin
      _T_4831_16 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_16 <= _T_4006_16;
      end
    end
    if (_T_337) begin
      _T_4831_17 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_17 <= _T_4006_17;
      end
    end
    if (_T_337) begin
      _T_4831_18 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_18 <= _T_4006_18;
      end
    end
    if (_T_337) begin
      _T_4831_19 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_19 <= _T_4006_19;
      end
    end
    if (_T_337) begin
      _T_4831_20 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_20 <= _T_4006_20;
      end
    end
    if (_T_337) begin
      _T_4831_21 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_21 <= _T_4006_21;
      end
    end
    if (_T_337) begin
      _T_4831_22 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_22 <= _T_4006_22;
      end
    end
    if (_T_337) begin
      _T_4831_23 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_23 <= _T_4006_23;
      end
    end
    if (_T_337) begin
      _T_4831_24 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_24 <= _T_4006_24;
      end
    end
    if (_T_337) begin
      _T_4831_25 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_25 <= _T_4006_25;
      end
    end
    if (_T_337) begin
      _T_4831_26 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_26 <= _T_4006_26;
      end
    end
    if (_T_337) begin
      _T_4831_27 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_27 <= _T_4006_27;
      end
    end
    if (_T_337) begin
      _T_4831_28 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_28 <= _T_4006_28;
      end
    end
    if (_T_337) begin
      _T_4831_29 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_29 <= _T_4006_29;
      end
    end
    if (_T_337) begin
      _T_4831_30 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_30 <= _T_4006_30;
      end
    end
    if (_T_337) begin
      _T_4831_31 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_31 <= _T_4006_31;
      end
    end
    if (_T_337) begin
      _T_4831_32 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_32 <= _T_4006_32;
      end
    end
    if (_T_337) begin
      _T_4831_33 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_33 <= _T_4006_33;
      end
    end
    if (_T_337) begin
      _T_4831_34 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_34 <= _T_4006_34;
      end
    end
    if (_T_337) begin
      _T_4831_35 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_35 <= _T_4006_35;
      end
    end
    if (_T_337) begin
      _T_4831_36 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_36 <= _T_4006_36;
      end
    end
    if (_T_337) begin
      _T_4831_37 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_37 <= _T_4006_37;
      end
    end
    if (_T_337) begin
      _T_4831_38 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_38 <= _T_4006_38;
      end
    end
    if (_T_337) begin
      _T_4831_39 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_39 <= _T_4006_39;
      end
    end
    if (_T_337) begin
      _T_4831_40 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_40 <= _T_4006_40;
      end
    end
    if (_T_337) begin
      _T_4831_41 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_41 <= _T_4006_41;
      end
    end
    if (_T_337) begin
      _T_4831_42 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_42 <= _T_4006_42;
      end
    end
    if (_T_337) begin
      _T_4831_43 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_43 <= _T_4006_43;
      end
    end
    if (_T_337) begin
      _T_4831_44 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_44 <= _T_4006_44;
      end
    end
    if (_T_337) begin
      _T_4831_45 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_45 <= _T_4006_45;
      end
    end
    if (_T_337) begin
      _T_4831_46 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_46 <= _T_4006_46;
      end
    end
    if (_T_337) begin
      _T_4831_47 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_47 <= _T_4006_47;
      end
    end
    if (_T_337) begin
      _T_4831_48 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_48 <= _T_4006_48;
      end
    end
    if (_T_337) begin
      _T_4831_49 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_49 <= _T_4006_49;
      end
    end
    if (_T_337) begin
      _T_4831_50 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_50 <= _T_4006_50;
      end
    end
    if (_T_337) begin
      _T_4831_51 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_51 <= _T_4006_51;
      end
    end
    if (_T_337) begin
      _T_4831_52 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_52 <= _T_4006_52;
      end
    end
    if (_T_337) begin
      _T_4831_53 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_53 <= _T_4006_53;
      end
    end
    if (_T_337) begin
      _T_4831_54 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_54 <= _T_4006_54;
      end
    end
    if (_T_337) begin
      _T_4831_55 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_55 <= _T_4006_55;
      end
    end
    if (_T_337) begin
      _T_4831_56 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_56 <= _T_4006_56;
      end
    end
    if (_T_337) begin
      _T_4831_57 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_57 <= _T_4006_57;
      end
    end
    if (_T_337) begin
      _T_4831_58 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_58 <= _T_4006_58;
      end
    end
    if (_T_337) begin
      _T_4831_59 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_59 <= _T_4006_59;
      end
    end
    if (_T_337) begin
      _T_4831_60 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_60 <= _T_4006_60;
      end
    end
    if (_T_337) begin
      _T_4831_61 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_61 <= _T_4006_61;
      end
    end
    if (_T_337) begin
      _T_4831_62 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_62 <= _T_4006_62;
      end
    end
    if (_T_337) begin
      _T_4831_63 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_4831_63 <= _T_4006_63;
      end
    end
    if (_T_337) begin
      _T_5358_0 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_0 <= _T_4006_0;
      end
    end
    if (_T_337) begin
      _T_5358_1 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_1 <= _T_4006_1;
      end
    end
    if (_T_337) begin
      _T_5358_2 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_2 <= _T_4006_2;
      end
    end
    if (_T_337) begin
      _T_5358_3 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_3 <= _T_4006_3;
      end
    end
    if (_T_337) begin
      _T_5358_4 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_4 <= _T_4006_4;
      end
    end
    if (_T_337) begin
      _T_5358_5 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_5 <= _T_4006_5;
      end
    end
    if (_T_337) begin
      _T_5358_6 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_6 <= _T_4006_6;
      end
    end
    if (_T_337) begin
      _T_5358_7 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_7 <= _T_4006_7;
      end
    end
    if (_T_337) begin
      _T_5358_8 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_8 <= _T_4006_8;
      end
    end
    if (_T_337) begin
      _T_5358_9 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_9 <= _T_4006_9;
      end
    end
    if (_T_337) begin
      _T_5358_10 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_10 <= _T_4006_10;
      end
    end
    if (_T_337) begin
      _T_5358_11 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_11 <= _T_4006_11;
      end
    end
    if (_T_337) begin
      _T_5358_12 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_12 <= _T_4006_12;
      end
    end
    if (_T_337) begin
      _T_5358_13 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_13 <= _T_4006_13;
      end
    end
    if (_T_337) begin
      _T_5358_14 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_14 <= _T_4006_14;
      end
    end
    if (_T_337) begin
      _T_5358_15 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_15 <= _T_4006_15;
      end
    end
    if (_T_337) begin
      _T_5358_16 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_16 <= _T_4006_16;
      end
    end
    if (_T_337) begin
      _T_5358_17 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_17 <= _T_4006_17;
      end
    end
    if (_T_337) begin
      _T_5358_18 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_18 <= _T_4006_18;
      end
    end
    if (_T_337) begin
      _T_5358_19 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_19 <= _T_4006_19;
      end
    end
    if (_T_337) begin
      _T_5358_20 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_20 <= _T_4006_20;
      end
    end
    if (_T_337) begin
      _T_5358_21 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_21 <= _T_4006_21;
      end
    end
    if (_T_337) begin
      _T_5358_22 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_22 <= _T_4006_22;
      end
    end
    if (_T_337) begin
      _T_5358_23 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_23 <= _T_4006_23;
      end
    end
    if (_T_337) begin
      _T_5358_24 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_24 <= _T_4006_24;
      end
    end
    if (_T_337) begin
      _T_5358_25 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_25 <= _T_4006_25;
      end
    end
    if (_T_337) begin
      _T_5358_26 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_26 <= _T_4006_26;
      end
    end
    if (_T_337) begin
      _T_5358_27 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_27 <= _T_4006_27;
      end
    end
    if (_T_337) begin
      _T_5358_28 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_28 <= _T_4006_28;
      end
    end
    if (_T_337) begin
      _T_5358_29 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_29 <= _T_4006_29;
      end
    end
    if (_T_337) begin
      _T_5358_30 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_30 <= _T_4006_30;
      end
    end
    if (_T_337) begin
      _T_5358_31 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_31 <= _T_4006_31;
      end
    end
    if (_T_337) begin
      _T_5358_32 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_32 <= _T_4006_32;
      end
    end
    if (_T_337) begin
      _T_5358_33 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_33 <= _T_4006_33;
      end
    end
    if (_T_337) begin
      _T_5358_34 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_34 <= _T_4006_34;
      end
    end
    if (_T_337) begin
      _T_5358_35 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_35 <= _T_4006_35;
      end
    end
    if (_T_337) begin
      _T_5358_36 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_36 <= _T_4006_36;
      end
    end
    if (_T_337) begin
      _T_5358_37 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_37 <= _T_4006_37;
      end
    end
    if (_T_337) begin
      _T_5358_38 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_38 <= _T_4006_38;
      end
    end
    if (_T_337) begin
      _T_5358_39 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_39 <= _T_4006_39;
      end
    end
    if (_T_337) begin
      _T_5358_40 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_40 <= _T_4006_40;
      end
    end
    if (_T_337) begin
      _T_5358_41 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_41 <= _T_4006_41;
      end
    end
    if (_T_337) begin
      _T_5358_42 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_42 <= _T_4006_42;
      end
    end
    if (_T_337) begin
      _T_5358_43 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_43 <= _T_4006_43;
      end
    end
    if (_T_337) begin
      _T_5358_44 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_44 <= _T_4006_44;
      end
    end
    if (_T_337) begin
      _T_5358_45 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_45 <= _T_4006_45;
      end
    end
    if (_T_337) begin
      _T_5358_46 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_46 <= _T_4006_46;
      end
    end
    if (_T_337) begin
      _T_5358_47 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_47 <= _T_4006_47;
      end
    end
    if (_T_337) begin
      _T_5358_48 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_48 <= _T_4006_48;
      end
    end
    if (_T_337) begin
      _T_5358_49 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_49 <= _T_4006_49;
      end
    end
    if (_T_337) begin
      _T_5358_50 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_50 <= _T_4006_50;
      end
    end
    if (_T_337) begin
      _T_5358_51 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_51 <= _T_4006_51;
      end
    end
    if (_T_337) begin
      _T_5358_52 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_52 <= _T_4006_52;
      end
    end
    if (_T_337) begin
      _T_5358_53 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_53 <= _T_4006_53;
      end
    end
    if (_T_337) begin
      _T_5358_54 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_54 <= _T_4006_54;
      end
    end
    if (_T_337) begin
      _T_5358_55 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_55 <= _T_4006_55;
      end
    end
    if (_T_337) begin
      _T_5358_56 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_56 <= _T_4006_56;
      end
    end
    if (_T_337) begin
      _T_5358_57 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_57 <= _T_4006_57;
      end
    end
    if (_T_337) begin
      _T_5358_58 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_58 <= _T_4006_58;
      end
    end
    if (_T_337) begin
      _T_5358_59 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_59 <= _T_4006_59;
      end
    end
    if (_T_337) begin
      _T_5358_60 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_60 <= _T_4006_60;
      end
    end
    if (_T_337) begin
      _T_5358_61 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_61 <= _T_4006_61;
      end
    end
    if (_T_337) begin
      _T_5358_62 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_62 <= _T_4006_62;
      end
    end
    if (_T_337) begin
      _T_5358_63 <= 1'h0;
    end else begin
      if (_T_4557) begin
        _T_5358_63 <= _T_4006_63;
      end
    end
    if (_T_4006_0) begin
      _T_5619 <= _T_4209_0;
    end
    if (_T_4006_0) begin
      _T_5621 <= _T_4209_0;
    end
    if (_T_4006_1) begin
      _T_5623 <= _T_4209_1;
    end
    if (_T_4006_1) begin
      _T_5625 <= _T_4209_1;
    end
    if (_T_4006_2) begin
      _T_5627 <= _T_4209_2;
    end
    if (_T_4006_2) begin
      _T_5629 <= _T_4209_2;
    end
    if (_T_4006_3) begin
      _T_5631 <= _T_4209_3;
    end
    if (_T_4006_3) begin
      _T_5633 <= _T_4209_3;
    end
    if (_T_4006_4) begin
      _T_5635 <= _T_4209_4;
    end
    if (_T_4006_4) begin
      _T_5637 <= _T_4209_4;
    end
    if (_T_4006_5) begin
      _T_5639 <= _T_4209_5;
    end
    if (_T_4006_5) begin
      _T_5641 <= _T_4209_5;
    end
    if (_T_4006_6) begin
      _T_5643 <= _T_4209_6;
    end
    if (_T_4006_6) begin
      _T_5645 <= _T_4209_6;
    end
    if (_T_4006_7) begin
      _T_5647 <= _T_4209_7;
    end
    if (_T_4006_7) begin
      _T_5649 <= _T_4209_7;
    end
    if (_T_4006_8) begin
      _T_5651 <= _T_4209_8;
    end
    if (_T_4006_8) begin
      _T_5653 <= _T_4209_8;
    end
    if (_T_4006_9) begin
      _T_5655 <= _T_4209_9;
    end
    if (_T_4006_9) begin
      _T_5657 <= _T_4209_9;
    end
    if (_T_4006_10) begin
      _T_5659 <= _T_4209_10;
    end
    if (_T_4006_10) begin
      _T_5661 <= _T_4209_10;
    end
    if (_T_4006_11) begin
      _T_5663 <= _T_4209_11;
    end
    if (_T_4006_11) begin
      _T_5665 <= _T_4209_11;
    end
    if (_T_4006_12) begin
      _T_5667 <= _T_4209_12;
    end
    if (_T_4006_12) begin
      _T_5669 <= _T_4209_12;
    end
    if (_T_4006_13) begin
      _T_5671 <= _T_4209_13;
    end
    if (_T_4006_13) begin
      _T_5673 <= _T_4209_13;
    end
    if (_T_4006_14) begin
      _T_5675 <= _T_4209_14;
    end
    if (_T_4006_14) begin
      _T_5677 <= _T_4209_14;
    end
    if (_T_4006_15) begin
      _T_5679 <= _T_4209_15;
    end
    if (_T_4006_15) begin
      _T_5681 <= _T_4209_15;
    end
    if (_T_4006_16) begin
      _T_5683 <= _T_4209_16;
    end
    if (_T_4006_16) begin
      _T_5685 <= _T_4209_16;
    end
    if (_T_4006_17) begin
      _T_5687 <= _T_4209_17;
    end
    if (_T_4006_17) begin
      _T_5689 <= _T_4209_17;
    end
    if (_T_4006_18) begin
      _T_5691 <= _T_4209_18;
    end
    if (_T_4006_18) begin
      _T_5693 <= _T_4209_18;
    end
    if (_T_4006_19) begin
      _T_5695 <= _T_4209_19;
    end
    if (_T_4006_19) begin
      _T_5697 <= _T_4209_19;
    end
    if (_T_4006_20) begin
      _T_5699 <= _T_4209_20;
    end
    if (_T_4006_20) begin
      _T_5701 <= _T_4209_20;
    end
    if (_T_4006_21) begin
      _T_5703 <= _T_4209_21;
    end
    if (_T_4006_21) begin
      _T_5705 <= _T_4209_21;
    end
    if (_T_4006_22) begin
      _T_5707 <= _T_4209_22;
    end
    if (_T_4006_22) begin
      _T_5709 <= _T_4209_22;
    end
    if (_T_4006_23) begin
      _T_5711 <= _T_4209_23;
    end
    if (_T_4006_23) begin
      _T_5713 <= _T_4209_23;
    end
    if (_T_4006_24) begin
      _T_5715 <= _T_4209_24;
    end
    if (_T_4006_24) begin
      _T_5717 <= _T_4209_24;
    end
    if (_T_4006_25) begin
      _T_5719 <= _T_4209_25;
    end
    if (_T_4006_25) begin
      _T_5721 <= _T_4209_25;
    end
    if (_T_4006_26) begin
      _T_5723 <= _T_4209_26;
    end
    if (_T_4006_26) begin
      _T_5725 <= _T_4209_26;
    end
    if (_T_4006_27) begin
      _T_5727 <= _T_4209_27;
    end
    if (_T_4006_27) begin
      _T_5729 <= _T_4209_27;
    end
    if (_T_4006_28) begin
      _T_5731 <= _T_4209_28;
    end
    if (_T_4006_28) begin
      _T_5733 <= _T_4209_28;
    end
    if (_T_4006_29) begin
      _T_5735 <= _T_4209_29;
    end
    if (_T_4006_29) begin
      _T_5737 <= _T_4209_29;
    end
    if (_T_4006_30) begin
      _T_5739 <= _T_4209_30;
    end
    if (_T_4006_30) begin
      _T_5741 <= _T_4209_30;
    end
    if (_T_4006_31) begin
      _T_5743 <= _T_4209_31;
    end
    if (_T_4006_31) begin
      _T_5745 <= _T_4209_31;
    end
    if (_T_4006_32) begin
      _T_5747 <= _T_4209_32;
    end
    if (_T_4006_32) begin
      _T_5749 <= _T_4209_32;
    end
    if (_T_4006_33) begin
      _T_5751 <= _T_4209_33;
    end
    if (_T_4006_33) begin
      _T_5753 <= _T_4209_33;
    end
    if (_T_4006_34) begin
      _T_5755 <= _T_4209_34;
    end
    if (_T_4006_34) begin
      _T_5757 <= _T_4209_34;
    end
    if (_T_4006_35) begin
      _T_5759 <= _T_4209_35;
    end
    if (_T_4006_35) begin
      _T_5761 <= _T_4209_35;
    end
    if (_T_4006_36) begin
      _T_5763 <= _T_4209_36;
    end
    if (_T_4006_36) begin
      _T_5765 <= _T_4209_36;
    end
    if (_T_4006_37) begin
      _T_5767 <= _T_4209_37;
    end
    if (_T_4006_37) begin
      _T_5769 <= _T_4209_37;
    end
    if (_T_4006_38) begin
      _T_5771 <= _T_4209_38;
    end
    if (_T_4006_38) begin
      _T_5773 <= _T_4209_38;
    end
    if (_T_4006_39) begin
      _T_5775 <= _T_4209_39;
    end
    if (_T_4006_39) begin
      _T_5777 <= _T_4209_39;
    end
    if (_T_4006_40) begin
      _T_5779 <= _T_4209_40;
    end
    if (_T_4006_40) begin
      _T_5781 <= _T_4209_40;
    end
    if (_T_4006_41) begin
      _T_5783 <= _T_4209_41;
    end
    if (_T_4006_41) begin
      _T_5785 <= _T_4209_41;
    end
    if (_T_4006_42) begin
      _T_5787 <= _T_4209_42;
    end
    if (_T_4006_42) begin
      _T_5789 <= _T_4209_42;
    end
    if (_T_4006_43) begin
      _T_5791 <= _T_4209_43;
    end
    if (_T_4006_43) begin
      _T_5793 <= _T_4209_43;
    end
    if (_T_4006_44) begin
      _T_5795 <= _T_4209_44;
    end
    if (_T_4006_44) begin
      _T_5797 <= _T_4209_44;
    end
    if (_T_4006_45) begin
      _T_5799 <= _T_4209_45;
    end
    if (_T_4006_45) begin
      _T_5801 <= _T_4209_45;
    end
    if (_T_4006_46) begin
      _T_5803 <= _T_4209_46;
    end
    if (_T_4006_46) begin
      _T_5805 <= _T_4209_46;
    end
    if (_T_4006_47) begin
      _T_5807 <= _T_4209_47;
    end
    if (_T_4006_47) begin
      _T_5809 <= _T_4209_47;
    end
    if (_T_4006_48) begin
      _T_5811 <= _T_4209_48;
    end
    if (_T_4006_48) begin
      _T_5813 <= _T_4209_48;
    end
    if (_T_4006_49) begin
      _T_5815 <= _T_4209_49;
    end
    if (_T_4006_49) begin
      _T_5817 <= _T_4209_49;
    end
    if (_T_4006_50) begin
      _T_5819 <= _T_4209_50;
    end
    if (_T_4006_50) begin
      _T_5821 <= _T_4209_50;
    end
    if (_T_4006_51) begin
      _T_5823 <= _T_4209_51;
    end
    if (_T_4006_51) begin
      _T_5825 <= _T_4209_51;
    end
    if (_T_4006_52) begin
      _T_5827 <= _T_4209_52;
    end
    if (_T_4006_52) begin
      _T_5829 <= _T_4209_52;
    end
    if (_T_4006_53) begin
      _T_5831 <= _T_4209_53;
    end
    if (_T_4006_53) begin
      _T_5833 <= _T_4209_53;
    end
    if (_T_4006_54) begin
      _T_5835 <= _T_4209_54;
    end
    if (_T_4006_54) begin
      _T_5837 <= _T_4209_54;
    end
    if (_T_4006_55) begin
      _T_5839 <= _T_4209_55;
    end
    if (_T_4006_55) begin
      _T_5841 <= _T_4209_55;
    end
    if (_T_4006_56) begin
      _T_5843 <= _T_4209_56;
    end
    if (_T_4006_56) begin
      _T_5845 <= _T_4209_56;
    end
    if (_T_4006_57) begin
      _T_5847 <= _T_4209_57;
    end
    if (_T_4006_57) begin
      _T_5849 <= _T_4209_57;
    end
    if (_T_4006_58) begin
      _T_5851 <= _T_4209_58;
    end
    if (_T_4006_58) begin
      _T_5853 <= _T_4209_58;
    end
    if (_T_4006_59) begin
      _T_5855 <= _T_4209_59;
    end
    if (_T_4006_59) begin
      _T_5857 <= _T_4209_59;
    end
    if (_T_4006_60) begin
      _T_5859 <= _T_4209_60;
    end
    if (_T_4006_60) begin
      _T_5861 <= _T_4209_60;
    end
    if (_T_4006_61) begin
      _T_5863 <= _T_4209_61;
    end
    if (_T_4006_61) begin
      _T_5865 <= _T_4209_61;
    end
    if (_T_4006_62) begin
      _T_5867 <= _T_4209_62;
    end
    if (_T_4006_62) begin
      _T_5869 <= _T_4209_62;
    end
    if (_T_4006_63) begin
      _T_5871 <= _T_4209_63;
    end
    if (_T_4006_63) begin
      _T_5873 <= _T_4209_63;
    end
  end
  always @(posedge nvdla_core_ng_clk) begin
    if (_T_337) begin
      _T_793 <= 15'h0;
    end else begin
      if (_T_865) begin
        if (sc2cdma_dat_pending_req) begin
          _T_793 <= 15'h0;
        end else begin
          if (_T_836) begin
            _T_793 <= _T_829;
          end else begin
            _T_793 <= _T_820;
          end
        end
      end
    end
  end
endmodule


// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CSC_dl.v
// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CSC.h

module NV_NVDLA_CSC_dl (
   nvdla_core_clk //|< i
  ,nvdla_core_rstn //|< i
  ,sg2dl_pvld //|< i
  ,sg2dl_pd //|< i
  ,sc_state //|< i
  ,sg2dl_reuse_rls //|< i
  ,sc2cdma_dat_pending_req //|< i
  ,cdma2sc_dat_updt //|< i
  ,cdma2sc_dat_entries //|< i
  ,cdma2sc_dat_slices //|< i
  ,sc2cdma_dat_updt //|> o
  ,sc2cdma_dat_entries //|> o
  ,sc2cdma_dat_slices //|> o
  ,sc2buf_dat_rd_en //|> o
  ,sc2buf_dat_rd_addr //|> o
  ,sc2buf_dat_rd_valid //|< i
  ,sc2buf_dat_rd_data //|< i
  ,sc2mac_dat_a_pvld //|> o
  ,sc2mac_dat_a_mask //|> o
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: ,sc2mac_dat_a_data${i} //|> o )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,sc2mac_dat_a_data0 //|> o 
,sc2mac_dat_a_data1 //|> o 
,sc2mac_dat_a_data2 //|> o 
,sc2mac_dat_a_data3 //|> o 
,sc2mac_dat_a_data4 //|> o 
,sc2mac_dat_a_data5 //|> o 
,sc2mac_dat_a_data6 //|> o 
,sc2mac_dat_a_data7 //|> o 
,sc2mac_dat_a_data8 //|> o 
,sc2mac_dat_a_data9 //|> o 
,sc2mac_dat_a_data10 //|> o 
,sc2mac_dat_a_data11 //|> o 
,sc2mac_dat_a_data12 //|> o 
,sc2mac_dat_a_data13 //|> o 
,sc2mac_dat_a_data14 //|> o 
,sc2mac_dat_a_data15 //|> o 
,sc2mac_dat_a_data16 //|> o 
,sc2mac_dat_a_data17 //|> o 
,sc2mac_dat_a_data18 //|> o 
,sc2mac_dat_a_data19 //|> o 
,sc2mac_dat_a_data20 //|> o 
,sc2mac_dat_a_data21 //|> o 
,sc2mac_dat_a_data22 //|> o 
,sc2mac_dat_a_data23 //|> o 
,sc2mac_dat_a_data24 //|> o 
,sc2mac_dat_a_data25 //|> o 
,sc2mac_dat_a_data26 //|> o 
,sc2mac_dat_a_data27 //|> o 
,sc2mac_dat_a_data28 //|> o 
,sc2mac_dat_a_data29 //|> o 
,sc2mac_dat_a_data30 //|> o 
,sc2mac_dat_a_data31 //|> o 
,sc2mac_dat_a_data32 //|> o 
,sc2mac_dat_a_data33 //|> o 
,sc2mac_dat_a_data34 //|> o 
,sc2mac_dat_a_data35 //|> o 
,sc2mac_dat_a_data36 //|> o 
,sc2mac_dat_a_data37 //|> o 
,sc2mac_dat_a_data38 //|> o 
,sc2mac_dat_a_data39 //|> o 
,sc2mac_dat_a_data40 //|> o 
,sc2mac_dat_a_data41 //|> o 
,sc2mac_dat_a_data42 //|> o 
,sc2mac_dat_a_data43 //|> o 
,sc2mac_dat_a_data44 //|> o 
,sc2mac_dat_a_data45 //|> o 
,sc2mac_dat_a_data46 //|> o 
,sc2mac_dat_a_data47 //|> o 
,sc2mac_dat_a_data48 //|> o 
,sc2mac_dat_a_data49 //|> o 
,sc2mac_dat_a_data50 //|> o 
,sc2mac_dat_a_data51 //|> o 
,sc2mac_dat_a_data52 //|> o 
,sc2mac_dat_a_data53 //|> o 
,sc2mac_dat_a_data54 //|> o 
,sc2mac_dat_a_data55 //|> o 
,sc2mac_dat_a_data56 //|> o 
,sc2mac_dat_a_data57 //|> o 
,sc2mac_dat_a_data58 //|> o 
,sc2mac_dat_a_data59 //|> o 
,sc2mac_dat_a_data60 //|> o 
,sc2mac_dat_a_data61 //|> o 
,sc2mac_dat_a_data62 //|> o 
,sc2mac_dat_a_data63 //|> o 
//| eperl: generated_end (DO NOT EDIT ABOVE)
  ,sc2mac_dat_a_pd //|> o
  ,sc2mac_dat_b_pvld //|> o
  ,sc2mac_dat_b_mask //|> o
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: ,sc2mac_dat_b_data${i} //|> o )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,sc2mac_dat_b_data0 //|> o 
,sc2mac_dat_b_data1 //|> o 
,sc2mac_dat_b_data2 //|> o 
,sc2mac_dat_b_data3 //|> o 
,sc2mac_dat_b_data4 //|> o 
,sc2mac_dat_b_data5 //|> o 
,sc2mac_dat_b_data6 //|> o 
,sc2mac_dat_b_data7 //|> o 
,sc2mac_dat_b_data8 //|> o 
,sc2mac_dat_b_data9 //|> o 
,sc2mac_dat_b_data10 //|> o 
,sc2mac_dat_b_data11 //|> o 
,sc2mac_dat_b_data12 //|> o 
,sc2mac_dat_b_data13 //|> o 
,sc2mac_dat_b_data14 //|> o 
,sc2mac_dat_b_data15 //|> o 
,sc2mac_dat_b_data16 //|> o 
,sc2mac_dat_b_data17 //|> o 
,sc2mac_dat_b_data18 //|> o 
,sc2mac_dat_b_data19 //|> o 
,sc2mac_dat_b_data20 //|> o 
,sc2mac_dat_b_data21 //|> o 
,sc2mac_dat_b_data22 //|> o 
,sc2mac_dat_b_data23 //|> o 
,sc2mac_dat_b_data24 //|> o 
,sc2mac_dat_b_data25 //|> o 
,sc2mac_dat_b_data26 //|> o 
,sc2mac_dat_b_data27 //|> o 
,sc2mac_dat_b_data28 //|> o 
,sc2mac_dat_b_data29 //|> o 
,sc2mac_dat_b_data30 //|> o 
,sc2mac_dat_b_data31 //|> o 
,sc2mac_dat_b_data32 //|> o 
,sc2mac_dat_b_data33 //|> o 
,sc2mac_dat_b_data34 //|> o 
,sc2mac_dat_b_data35 //|> o 
,sc2mac_dat_b_data36 //|> o 
,sc2mac_dat_b_data37 //|> o 
,sc2mac_dat_b_data38 //|> o 
,sc2mac_dat_b_data39 //|> o 
,sc2mac_dat_b_data40 //|> o 
,sc2mac_dat_b_data41 //|> o 
,sc2mac_dat_b_data42 //|> o 
,sc2mac_dat_b_data43 //|> o 
,sc2mac_dat_b_data44 //|> o 
,sc2mac_dat_b_data45 //|> o 
,sc2mac_dat_b_data46 //|> o 
,sc2mac_dat_b_data47 //|> o 
,sc2mac_dat_b_data48 //|> o 
,sc2mac_dat_b_data49 //|> o 
,sc2mac_dat_b_data50 //|> o 
,sc2mac_dat_b_data51 //|> o 
,sc2mac_dat_b_data52 //|> o 
,sc2mac_dat_b_data53 //|> o 
,sc2mac_dat_b_data54 //|> o 
,sc2mac_dat_b_data55 //|> o 
,sc2mac_dat_b_data56 //|> o 
,sc2mac_dat_b_data57 //|> o 
,sc2mac_dat_b_data58 //|> o 
,sc2mac_dat_b_data59 //|> o 
,sc2mac_dat_b_data60 //|> o 
,sc2mac_dat_b_data61 //|> o 
,sc2mac_dat_b_data62 //|> o 
,sc2mac_dat_b_data63 //|> o 
//| eperl: generated_end (DO NOT EDIT ABOVE)
  ,sc2mac_dat_b_pd //|> o
  ,nvdla_core_ng_clk //|< i
  ,reg2dp_op_en //|< i
  ,reg2dp_conv_mode //|< i
  ,reg2dp_batches //|< i
  ,reg2dp_proc_precision //|< i
  ,reg2dp_datain_format //|< i
  ,reg2dp_skip_data_rls //|< i
  ,reg2dp_datain_channel_ext //|< i
  ,reg2dp_datain_height_ext //|< i
  ,reg2dp_datain_width_ext //|< i
  ,reg2dp_y_extension //|< i
  ,reg2dp_weight_channel_ext //|< i
  ,reg2dp_entries //|< i
  ,reg2dp_dataout_width //|< i
  ,reg2dp_rls_slices //|< i
  ,reg2dp_conv_x_stride_ext //|< i
  ,reg2dp_conv_y_stride_ext //|< i
  ,reg2dp_x_dilation_ext //|< i
  ,reg2dp_y_dilation_ext //|< i
  ,reg2dp_pad_left //|< i
  ,reg2dp_pad_top //|< i
  ,reg2dp_pad_value //|< i
  ,reg2dp_data_bank //|< i
  ,reg2dp_pra_truncate //|< i
  ,slcg_wg_en //|> o
  );
input nvdla_core_clk;
input nvdla_core_rstn;
input sg2dl_pvld; /* data valid */
input [30:0] sg2dl_pd;
input [1:0] sc_state;
input sg2dl_reuse_rls;
input sc2cdma_dat_pending_req;
input cdma2sc_dat_updt; /* data valid */
input [15 -1:0] cdma2sc_dat_entries;
input [13:0] cdma2sc_dat_slices;
output sc2cdma_dat_updt; /* data valid */
output [15 -1:0] sc2cdma_dat_entries;
output [13:0] sc2cdma_dat_slices;
output sc2buf_dat_rd_en; /* data valid */
output [13 -1:0] sc2buf_dat_rd_addr;
input sc2buf_dat_rd_valid; /* data valid */
input [512 -1:0] sc2buf_dat_rd_data;
output sc2mac_dat_a_pvld; /* data valid */
output [64 -1:0] sc2mac_dat_a_mask;
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: output [8 -1:0] sc2mac_dat_a_data${i}; )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

output [8 -1:0] sc2mac_dat_a_data0; 
output [8 -1:0] sc2mac_dat_a_data1; 
output [8 -1:0] sc2mac_dat_a_data2; 
output [8 -1:0] sc2mac_dat_a_data3; 
output [8 -1:0] sc2mac_dat_a_data4; 
output [8 -1:0] sc2mac_dat_a_data5; 
output [8 -1:0] sc2mac_dat_a_data6; 
output [8 -1:0] sc2mac_dat_a_data7; 
output [8 -1:0] sc2mac_dat_a_data8; 
output [8 -1:0] sc2mac_dat_a_data9; 
output [8 -1:0] sc2mac_dat_a_data10; 
output [8 -1:0] sc2mac_dat_a_data11; 
output [8 -1:0] sc2mac_dat_a_data12; 
output [8 -1:0] sc2mac_dat_a_data13; 
output [8 -1:0] sc2mac_dat_a_data14; 
output [8 -1:0] sc2mac_dat_a_data15; 
output [8 -1:0] sc2mac_dat_a_data16; 
output [8 -1:0] sc2mac_dat_a_data17; 
output [8 -1:0] sc2mac_dat_a_data18; 
output [8 -1:0] sc2mac_dat_a_data19; 
output [8 -1:0] sc2mac_dat_a_data20; 
output [8 -1:0] sc2mac_dat_a_data21; 
output [8 -1:0] sc2mac_dat_a_data22; 
output [8 -1:0] sc2mac_dat_a_data23; 
output [8 -1:0] sc2mac_dat_a_data24; 
output [8 -1:0] sc2mac_dat_a_data25; 
output [8 -1:0] sc2mac_dat_a_data26; 
output [8 -1:0] sc2mac_dat_a_data27; 
output [8 -1:0] sc2mac_dat_a_data28; 
output [8 -1:0] sc2mac_dat_a_data29; 
output [8 -1:0] sc2mac_dat_a_data30; 
output [8 -1:0] sc2mac_dat_a_data31; 
output [8 -1:0] sc2mac_dat_a_data32; 
output [8 -1:0] sc2mac_dat_a_data33; 
output [8 -1:0] sc2mac_dat_a_data34; 
output [8 -1:0] sc2mac_dat_a_data35; 
output [8 -1:0] sc2mac_dat_a_data36; 
output [8 -1:0] sc2mac_dat_a_data37; 
output [8 -1:0] sc2mac_dat_a_data38; 
output [8 -1:0] sc2mac_dat_a_data39; 
output [8 -1:0] sc2mac_dat_a_data40; 
output [8 -1:0] sc2mac_dat_a_data41; 
output [8 -1:0] sc2mac_dat_a_data42; 
output [8 -1:0] sc2mac_dat_a_data43; 
output [8 -1:0] sc2mac_dat_a_data44; 
output [8 -1:0] sc2mac_dat_a_data45; 
output [8 -1:0] sc2mac_dat_a_data46; 
output [8 -1:0] sc2mac_dat_a_data47; 
output [8 -1:0] sc2mac_dat_a_data48; 
output [8 -1:0] sc2mac_dat_a_data49; 
output [8 -1:0] sc2mac_dat_a_data50; 
output [8 -1:0] sc2mac_dat_a_data51; 
output [8 -1:0] sc2mac_dat_a_data52; 
output [8 -1:0] sc2mac_dat_a_data53; 
output [8 -1:0] sc2mac_dat_a_data54; 
output [8 -1:0] sc2mac_dat_a_data55; 
output [8 -1:0] sc2mac_dat_a_data56; 
output [8 -1:0] sc2mac_dat_a_data57; 
output [8 -1:0] sc2mac_dat_a_data58; 
output [8 -1:0] sc2mac_dat_a_data59; 
output [8 -1:0] sc2mac_dat_a_data60; 
output [8 -1:0] sc2mac_dat_a_data61; 
output [8 -1:0] sc2mac_dat_a_data62; 
output [8 -1:0] sc2mac_dat_a_data63; 
//| eperl: generated_end (DO NOT EDIT ABOVE)
output [8:0] sc2mac_dat_a_pd;
output sc2mac_dat_b_pvld; /* data valid */
output [64 -1:0] sc2mac_dat_b_mask;
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: output [8 -1:0] sc2mac_dat_b_data${i}; )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

output [8 -1:0] sc2mac_dat_b_data0; 
output [8 -1:0] sc2mac_dat_b_data1; 
output [8 -1:0] sc2mac_dat_b_data2; 
output [8 -1:0] sc2mac_dat_b_data3; 
output [8 -1:0] sc2mac_dat_b_data4; 
output [8 -1:0] sc2mac_dat_b_data5; 
output [8 -1:0] sc2mac_dat_b_data6; 
output [8 -1:0] sc2mac_dat_b_data7; 
output [8 -1:0] sc2mac_dat_b_data8; 
output [8 -1:0] sc2mac_dat_b_data9; 
output [8 -1:0] sc2mac_dat_b_data10; 
output [8 -1:0] sc2mac_dat_b_data11; 
output [8 -1:0] sc2mac_dat_b_data12; 
output [8 -1:0] sc2mac_dat_b_data13; 
output [8 -1:0] sc2mac_dat_b_data14; 
output [8 -1:0] sc2mac_dat_b_data15; 
output [8 -1:0] sc2mac_dat_b_data16; 
output [8 -1:0] sc2mac_dat_b_data17; 
output [8 -1:0] sc2mac_dat_b_data18; 
output [8 -1:0] sc2mac_dat_b_data19; 
output [8 -1:0] sc2mac_dat_b_data20; 
output [8 -1:0] sc2mac_dat_b_data21; 
output [8 -1:0] sc2mac_dat_b_data22; 
output [8 -1:0] sc2mac_dat_b_data23; 
output [8 -1:0] sc2mac_dat_b_data24; 
output [8 -1:0] sc2mac_dat_b_data25; 
output [8 -1:0] sc2mac_dat_b_data26; 
output [8 -1:0] sc2mac_dat_b_data27; 
output [8 -1:0] sc2mac_dat_b_data28; 
output [8 -1:0] sc2mac_dat_b_data29; 
output [8 -1:0] sc2mac_dat_b_data30; 
output [8 -1:0] sc2mac_dat_b_data31; 
output [8 -1:0] sc2mac_dat_b_data32; 
output [8 -1:0] sc2mac_dat_b_data33; 
output [8 -1:0] sc2mac_dat_b_data34; 
output [8 -1:0] sc2mac_dat_b_data35; 
output [8 -1:0] sc2mac_dat_b_data36; 
output [8 -1:0] sc2mac_dat_b_data37; 
output [8 -1:0] sc2mac_dat_b_data38; 
output [8 -1:0] sc2mac_dat_b_data39; 
output [8 -1:0] sc2mac_dat_b_data40; 
output [8 -1:0] sc2mac_dat_b_data41; 
output [8 -1:0] sc2mac_dat_b_data42; 
output [8 -1:0] sc2mac_dat_b_data43; 
output [8 -1:0] sc2mac_dat_b_data44; 
output [8 -1:0] sc2mac_dat_b_data45; 
output [8 -1:0] sc2mac_dat_b_data46; 
output [8 -1:0] sc2mac_dat_b_data47; 
output [8 -1:0] sc2mac_dat_b_data48; 
output [8 -1:0] sc2mac_dat_b_data49; 
output [8 -1:0] sc2mac_dat_b_data50; 
output [8 -1:0] sc2mac_dat_b_data51; 
output [8 -1:0] sc2mac_dat_b_data52; 
output [8 -1:0] sc2mac_dat_b_data53; 
output [8 -1:0] sc2mac_dat_b_data54; 
output [8 -1:0] sc2mac_dat_b_data55; 
output [8 -1:0] sc2mac_dat_b_data56; 
output [8 -1:0] sc2mac_dat_b_data57; 
output [8 -1:0] sc2mac_dat_b_data58; 
output [8 -1:0] sc2mac_dat_b_data59; 
output [8 -1:0] sc2mac_dat_b_data60; 
output [8 -1:0] sc2mac_dat_b_data61; 
output [8 -1:0] sc2mac_dat_b_data62; 
output [8 -1:0] sc2mac_dat_b_data63; 
//| eperl: generated_end (DO NOT EDIT ABOVE)
output [8:0] sc2mac_dat_b_pd;
input nvdla_core_ng_clk;
input [0:0] reg2dp_op_en;
input [0:0] reg2dp_conv_mode;
input [4:0] reg2dp_batches;
input [1:0] reg2dp_proc_precision;
input [0:0] reg2dp_datain_format;
input [0:0] reg2dp_skip_data_rls;
input [12:0] reg2dp_datain_channel_ext;
input [12:0] reg2dp_datain_height_ext;
input [12:0] reg2dp_datain_width_ext;
input [1:0] reg2dp_y_extension;
input [12:0] reg2dp_weight_channel_ext;
input [13:0] reg2dp_entries;
input [12:0] reg2dp_dataout_width;
input [11:0] reg2dp_rls_slices;
input [2:0] reg2dp_conv_x_stride_ext;
input [2:0] reg2dp_conv_y_stride_ext;
input [4:0] reg2dp_x_dilation_ext;
input [4:0] reg2dp_y_dilation_ext;
input [4:0] reg2dp_pad_left;
input [4:0] reg2dp_pad_top;
input [15:0] reg2dp_pad_value;
input [4:0] reg2dp_data_bank;
input [1:0] reg2dp_pra_truncate;
output slcg_wg_en;
reg [4:0] batch_cmp;
reg [4:0] batch_cnt;
reg [13 -1:0] c_bias;
reg [13 -1:0] c_bias_d1;
reg [3:0] conv_x_stride;
reg [3:0] conv_y_stride;
reg [15 -1:0] dat_entry_avl;
reg [15 -1:0] dat_entry_end;
reg [15 -1:0] dat_entry_st;
reg dat_exec_valid_d1;
reg dat_exec_valid_d2;
reg dat_l0c0_dummy;
reg [512 -1:0] dat_l0c0;
reg dat_l0c1_dummy;
reg [512 -1:0] dat_l0c1;
reg dat_l1c0_dummy;
reg [512 -1:0] dat_l1c0;
reg dat_l1c1_dummy;
reg [512 -1:0] dat_l1c1;
reg dat_l2c0_dummy;
reg [512 -1:0] dat_l2c0;
reg dat_l2c1_dummy;
reg [512 -1:0] dat_l2c1;
reg dat_l3c0_dummy;
reg [512 -1:0] dat_l3c0;
reg dat_l3c1_dummy;
reg [512 -1:0] dat_l3c1;
reg [512 -1:0] dat_out_bypass_data;
reg [64 -1:0] dat_out_bypass_mask;
reg [8:0] dat_out_flag;
reg dat_out_pvld;
reg dat_pipe_local_valid;
reg dat_pipe_valid_d1;
reg dat_pipe_valid_d2;
reg [7:0] dat_req_bytes_d1;
reg [7:0] dat_req_bytes_d2;
reg dat_req_ch_end_d1;
reg dat_req_ch_end_d2;
reg [1:0] dat_req_cur_sub_h_d1;
reg [1:0] dat_req_cur_sub_h_d2;
reg dat_req_dummy_d1;
reg dat_req_dummy_d2;
reg [8:0] dat_req_flag_d1;
reg [8:0] dat_req_flag_d2;
reg dat_req_rls_d1;
reg dat_req_rls_d2;
reg dat_req_sub_c_d1;
reg dat_req_sub_c_d2;
reg [13 -1:0] dat_req_sub_h_0_addr;
reg [13 -1:0] dat_req_sub_h_1_addr;
reg [13 -1:0] dat_req_sub_h_2_addr;
reg [13 -1:0] dat_req_sub_h_3_addr;
reg [1:0] dat_req_sub_h_d1;
reg [1:0] dat_req_sub_h_d2;
reg [1:0] dat_req_sub_w_d1;
reg [1:0] dat_req_sub_w_d2;
reg dat_req_sub_w_st_d1;
reg dat_req_sub_w_st_d2;
reg dat_req_valid_d1;
wire [512 -1:0] dat_rsp_l0_sft;
reg [512 -1:0] dat_rsp_l0_sft_d1;
reg [512 -1:0] dat_rsp_l0_sft_d2;
reg [512 -1:0] dat_rsp_l0_sft_d3;
wire [512 -1:0] dat_rsp_l1_sft;
reg [512 -1:0] dat_rsp_l1_sft_d2;
reg [512 -1:0] dat_rsp_l1_sft_d3;
wire [512 -1:0] dat_rsp_l2_sft;
reg [512 -1:0] dat_rsp_l2_sft_d3;
wire [512 -1:0] dat_rsp_l3_sft;
reg [26:0] dat_rsp_pd_d1;
reg [26:0] dat_rsp_pd_d2;
reg [26:0] dat_rsp_pd_d3;
reg [26:0] dat_rsp_pd_d4;
reg [3:0] dat_rsp_pra_en_d1;
reg dat_rsp_pvld_d1;
reg dat_rsp_pvld_d2;
reg dat_rsp_pvld_d3;
reg dat_rsp_pvld_d4;
reg [255:0] dat_rsp_wg_ch0_d1;
reg [255:0] dat_rsp_wg_ch1_d1;
reg [255:0] dat_rsp_wg_ch2_d1;
reg [255:0] dat_rsp_wg_ch3_d1;
reg [13:0] dat_slice_avl;
reg [4:0] data_bank;
reg [5:0] data_batch;
reg [10:0] datain_c_cnt;
reg [10:0] datain_channel_cmp;
reg [13:0] datain_h_cnt;
reg [13:0] datain_h_ori;
reg [12:0] datain_height_cmp;
reg [13:0] datain_w_cnt;
reg [13:0] datain_w_ori;
reg [13:0] datain_width;
reg [12:0] datain_width_cmp;
reg [12:0] dataout_w_cnt;
reg [12:0] dataout_w_ori;
reg [12:0] dataout_width_cmp;
reg [8:0] dl_out_flag;
reg [64 -1:0] dl_out_mask;
reg dl_out_pvld;
reg dl_out_pvld_d1;
reg [30:0] dl_pd_d1;
reg [30:0] dl_pd_d2;
reg [30:0] dl_pd_d3;
reg [30:0] dl_pd_d4;
reg dl_pvld_d1;
reg dl_pvld_d2;
reg dl_pvld_d3;
reg dl_pvld_d4;
reg [15 -1:0] entries;
reg [15 -1:0] entries_batch;
reg [15 -1:0] entries_cmp;
reg [13 -1:0] h_bias_0_d1;
reg [13 -1:0] h_bias_0_stride;
reg [13 -1:0] h_bias_1_d1;
reg [13 -1:0] h_bias_1_stride;
reg [13 -1:0] h_bias_2_d1;
reg [13 -1:0] h_bias_2_stride;
reg [13 -1:0] h_bias_3_d1;
reg [13 -1:0] h_bias_3_stride;
reg [13:0] h_offset_slice;
reg [33:0] is_img_d1;
reg is_sg_running_d1;
reg [21:0] is_winograd_d1;
reg [15 -1:0] last_entries;
reg [13:0] last_slices;
reg layer_st_d1;
reg [15:0] pad_value;
reg [11:0] pixel_ch_stride;
reg pixel_force_clr_d1;
reg pixel_force_fetch_d1;
reg [15:0] pixel_w_ch_ori;
reg [15:0] pixel_w_cnt;
reg [15:0] pixel_w_ori;
reg [6:0] pixel_x_add;
reg [6:0] pixel_x_byte_stride;
reg [5:0] pixel_x_init;
reg [6:0] pixel_x_init_offset;
reg pixel_x_stride_odd;
reg [7:0] pra_precision;
reg [7:0] pra_truncate;
reg [15 -1:0] rls_entries;
reg [13:0] rls_slices;
reg [7:0] rsp_sft_cnt_l0;
reg [7:0] rsp_sft_cnt_l0_ori;
reg [7:0] rsp_sft_cnt_l1;
reg [7:0] rsp_sft_cnt_l1_ori;
reg [7:0] rsp_sft_cnt_l2;
reg [7:0] rsp_sft_cnt_l2_ori;
reg [7:0] rsp_sft_cnt_l3;
reg [7:0] rsp_sft_cnt_l3_ori;
reg [13 -1:0] sc2buf_dat_rd_addr;
reg [13 -1:0] sc2buf_dat_rd_next1_addr;
reg sc2buf_dat_rd_en;
reg [15 -1:0] sc2cdma_dat_entries;
reg [13:0] sc2cdma_dat_slices;
reg sc2cdma_dat_updt;
reg [64 -1:0] sc2mac_dat_a_mask;
reg [8:0] sc2mac_dat_a_pd;
reg sc2mac_dat_a_pvld;
reg [64 -1:0] sc2mac_dat_b_mask;
reg [8:0] sc2mac_dat_b_pd;
reg sc2mac_dat_b_pvld;
reg slcg_wg_en_d1;
reg slcg_wg_en_d2;
reg slcg_wg_en_d3;
reg [13:0] slice_left;
reg [6:0] stripe_cnt;
reg [2:0] sub_h_cmp_g0;
reg [2:0] sub_h_cmp_g1;
reg [1:0] sub_h_cnt;
reg [2:0] sub_h_total_g0;
reg [2:0] sub_h_total_g1;
reg [2:0] sub_h_total_g10;
reg [2:0] sub_h_total_g11;
reg [1:0] sub_h_total_g2;
reg [2:0] sub_h_total_g3;
reg [2:0] sub_h_total_g4;
reg [2:0] sub_h_total_g5;
reg [2:0] sub_h_total_g6;
reg [2:0] sub_h_total_g7;
reg [2:0] sub_h_total_g8;
reg [2:0] sub_h_total_g9;
reg [13 -1:0] w_bias_d1;
reg [5:0] x_dilate;
reg [5:0] y_dilate;
wire [4:0] batch_cmp_w;
wire [4:0] batch_cnt_w;
wire [13 -1:0] c_bias_add;
wire c_bias_d1_reg_en;
wire c_bias_reg_en;
wire [13 -1:0] c_bias_w;
wire cbuf_reset;
wire [3:0] conv_x_stride_w;
wire [3:0] conv_y_stride_w;
wire dat_conv_req_dummy;
wire dat_dummy_l0_en;
wire dat_dummy_l1_en;
wire dat_dummy_l2_en;
wire dat_dummy_l3_en;
wire [15 -1:0] dat_entry_avl_add;
wire [15 -1:0] dat_entry_avl_sub;
wire [15 -1:0] dat_entry_avl_w;
wire [15 -1:0] dat_entry_end_inc;
wire [15 -1:0] dat_entry_end_inc_wrap;
wire [15 -1:0] dat_entry_end_w;
wire [15 -1:0] dat_entry_st_inc;
wire [15 -1:0] dat_entry_st_inc_wrap;
wire [15 -1:0] dat_entry_st_w;
wire mon_dat_entry_end_inc;
wire mon_dat_entry_st_inc;
wire dat_exec_valid;
wire dat_img_req_dummy;
wire dat_img_req_skip;
wire dat_l0_set;
wire dat_l0c0_dummy_w;
wire dat_l0c0_en;
wire dat_l0c1_dummy_w;
wire dat_l0c1_en;
wire dat_l1_set;
wire dat_l1c0_dummy_w;
wire dat_l1c0_en;
wire dat_l1c0_hi_en;
wire dat_l1c1_dummy_w;
wire dat_l1c1_en;
wire dat_l1c1_hi_en;
wire dat_l2_set;
wire dat_l2c0_dummy_w;
wire dat_l2c0_en;
wire dat_l2c1_dummy_w;
wire dat_l2c1_en;
wire dat_l3_set;
wire dat_l3c0_dummy_w;
wire dat_l3c0_en;
wire dat_l3c1_dummy_w;
wire dat_l3c1_en;
wire [512 -1:0] dat_out_bypass_data_w;
wire [64 -1:0] dat_out_bypass_mask_w;
wire dat_out_bypass_p0_vld_w;
wire [512 -1:0] dat_out_data;
wire [8:0] dat_out_flag_l0;
wire [8:0] dat_out_flag_w;
wire [64 -1:0] dat_out_mask;
wire dat_out_pvld_l0;
wire dat_out_pvld_w;
wire [512 -1:0] dat_out_wg_8b;
wire [512 -1:0] dat_out_wg_data;
wire [64 -1:0] dat_out_wg_mask;
wire [64 -1:0] dat_out_wg_mask_int8;
wire dat_pipe_local_valid_w;
wire dat_pipe_valid;
wire [512 -1:0] dat_pra_dat;
wire [255:0] dat_pra_dat_ch0;
wire [255:0] dat_pra_dat_ch1;
wire [255:0] dat_pra_dat_ch2;
wire [255:0] dat_pra_dat_ch3;
wire [13 -1:0] dat_req_addr_last;
wire [13:0] dat_req_addr_sum;
wire [13 -1:0] dat_req_addr_w;
wire [13 -1:0] dat_req_addr_wrap;
wire [13 -1:0] dat_req_base_d1;
wire mon_dat_req_addr_sum;
wire [4:0] dat_req_batch_index;
wire [7:0] dat_req_bytes;
wire dat_req_channel_end;
wire dat_req_dummy;
wire dat_req_exec_dummy;
wire dat_req_exec_pvld;
wire [1:0] dat_req_exec_sub_h;
wire [8:0] dat_req_flag_w;
wire dat_req_layer_end;
wire [7:0] dat_req_pipe_bytes;
wire dat_req_pipe_ch_end;
wire [1:0] dat_req_pipe_cur_sub_h;
wire dat_req_pipe_dummy;
wire [8:0] dat_req_pipe_flag;
wire [28:0] dat_req_pipe_pd;
wire dat_req_pipe_pvld;
wire dat_req_pipe_rls;
wire dat_req_pipe_sub_c;
wire [1:0] dat_req_pipe_sub_h;
wire [1:0] dat_req_pipe_sub_w;
wire dat_req_pipe_sub_w_st;
wire dat_req_skip;
wire dat_req_stripe_end;
wire dat_req_stripe_st;
wire dat_req_sub_c_w;
wire dat_req_sub_h_0_addr_en;
wire dat_req_sub_h_1_addr_en;
wire dat_req_sub_h_2_addr_en;
wire dat_req_sub_h_3_addr_en;
wire dat_req_sub_w_st_en;
wire [1:0] dat_req_sub_w_w;
wire dat_req_valid;
wire dat_rls;
wire [4:0] dat_rsp_batch_index;
wire [7:0] dat_rsp_bytes;
wire dat_rsp_ch_end;
wire dat_rsp_channel_end;
wire [512 -1:0] dat_rsp_conv;
wire [512 -1:0] dat_rsp_conv_8b;
wire [64 -1:0] dat_rsp_cur_h_e2_mask_8b;
wire [64 -1:0] dat_rsp_cur_h_e4_mask_8b;
wire [64 -1:0] dat_rsp_cur_h_mask_p1;
wire [31:0] dat_rsp_cur_h_mask_p2;
wire [31:0] dat_rsp_cur_h_mask_p3;
wire [1:0] dat_rsp_cur_sub_h;
wire [512 -1:0] dat_rsp_data_w;
wire dat_rsp_exec_dummy;
wire dat_rsp_exec_dummy_d0;
wire dat_rsp_exec_pvld;
wire dat_rsp_exec_pvld_d0;
wire [1:0] dat_rsp_exec_sub_h;
wire [1:0] dat_rsp_exec_sub_h_d0;
wire [8:0] dat_rsp_flag;
wire [512 -1:0] dat_rsp_img;
wire [512 -1:0] dat_rsp_img_8b;
wire dat_rsp_l0_block_end;
wire [8:0] dat_rsp_l0_flag;
wire dat_rsp_l0_pvld;
wire [512*2 -1:0] dat_rsp_l0_sft_in;
wire dat_rsp_l0_stripe_end;
wire dat_rsp_l0_sub_c;
wire [512 -1:0] dat_rsp_l0c0;
wire [512 -1:0] dat_rsp_l0c1;
wire dat_rsp_l1_block_end;
wire [8:0] dat_rsp_l1_flag;
wire dat_rsp_l1_pvld;
wire [512*2 -1:0] dat_rsp_l1_sft_in;
wire dat_rsp_l1_stripe_end;
wire dat_rsp_l1_sub_c;
wire [512 -1:0] dat_rsp_l1c0;
wire [512 -1:0] dat_rsp_l1c1;
wire dat_rsp_l2_block_end;
wire [8:0] dat_rsp_l2_flag;
wire dat_rsp_l2_pvld;
wire [512*2 -1:0] dat_rsp_l2_sft_in;
wire dat_rsp_l2_stripe_end;
wire dat_rsp_l2_sub_c;
wire [512 -1:0] dat_rsp_l2c0;
wire [512 -1:0] dat_rsp_l2c1;
wire dat_rsp_l3_block_end;
wire [8:0] dat_rsp_l3_flag;
wire dat_rsp_l3_pvld;
wire [512*2 -1:0] dat_rsp_l3_sft_in;
wire dat_rsp_l3_stripe_end;
wire dat_rsp_l3_sub_c;
wire [512 -1:0] dat_rsp_l3c0;
wire [512 -1:0] dat_rsp_l3c1;
wire dat_rsp_layer_end;
wire [64 -1:0] dat_rsp_mask_8b;
wire [64 -1:0] dat_rsp_mask_val_int8;
wire [64 -1:0] dat_rsp_mask_w;
wire [64 -1:0] dat_rsp_ori_mask;
wire dat_rsp_p0_vld_w;
wire dat_rsp_p1_vld_w;
wire [512 -1:0] dat_rsp_pad_value;
wire [26:0] dat_rsp_pd;
wire [26:0] dat_rsp_pd_d0;
wire [7:0] dat_rsp_pipe_bytes;
wire dat_rsp_pipe_ch_end;
wire [1:0] dat_rsp_pipe_cur_sub_h;
wire dat_rsp_pipe_dummy;
wire [8:0] dat_rsp_pipe_flag;
wire [28:0] dat_rsp_pipe_pd;
wire [28:0] dat_rsp_pipe_pd_d0;
wire dat_rsp_pipe_pvld;
wire dat_rsp_pipe_pvld_d0;
wire dat_rsp_pipe_rls;
wire dat_rsp_pipe_sub_c;
wire [1:0] dat_rsp_pipe_sub_h;
wire [1:0] dat_rsp_pipe_sub_w;
wire dat_rsp_pipe_sub_w_st;
wire dat_rsp_pra_en;
wire dat_rsp_pvld;
wire dat_rsp_pvld_d0;
wire dat_rsp_rls;
wire dat_rsp_stripe_end;
wire dat_rsp_stripe_st;
wire dat_rsp_sub_c;
wire [1:0] dat_rsp_sub_h;
wire [1:0] dat_rsp_sub_w;
wire [512 -1:0] dat_rsp_wg;
wire [255:0] dat_rsp_wg_ch0;
wire [255:0] dat_rsp_wg_ch1;
wire [255:0] dat_rsp_wg_ch2;
wire [255:0] dat_rsp_wg_ch3;
wire [512 -1:0] dat_rsp_wg_lb;
wire [512 -1:0] dat_rsp_wg_lt;
wire [512 -1:0] dat_rsp_wg_rb;
wire [512 -1:0] dat_rsp_wg_rt;
wire dat_rsp_wg_sel_8b_hi;
wire dat_rsp_wg_sel_8b_lo;
wire dat_rsp_wg_sel_lb;
wire dat_rsp_wg_sel_lt;
wire dat_rsp_wg_sel_rb;
wire dat_rsp_wg_sel_rt;
wire [13:0] dat_slice_avl_add;
wire [13:0] dat_slice_avl_sub;
wire [13:0] dat_slice_avl_w;
wire [2303:0] dat_wg;
wire [255:0] dat_wg_8b_ch0;
wire [255:0] dat_wg_8b_ch1;
wire [255:0] dat_wg_8b_ch2;
wire [255:0] dat_wg_8b_ch3;
wire [255:0] dat_wg_8b_ch4;
wire [255:0] dat_wg_8b_ch5;
wire [255:0] dat_wg_8b_ch6;
wire [255:0] dat_wg_8b_ch7;
wire dat_wg_adv;
wire dat_wg_req_dummy;
wire dat_wg_req_skip;
wire [4:0] data_bank_w;
wire [5:0] data_batch_w;
wire [10:0] datain_c_cnt_inc;
wire datain_c_cnt_reg_en;
wire [10:0] datain_c_cnt_w;
wire [10:0] datain_channel_cmp_w;
wire [13:0] datain_h_cnt_inc;
wire datain_h_cnt_reg_en;
wire [13:0] datain_h_cnt_st;
wire [13:0] datain_h_cnt_w;
wire [13:0] datain_h_cur;
wire datain_h_ori_reg_en;
wire [12:0] datain_height_cmp_w;
wire [13:0] datain_w_cnt_inc;
wire datain_w_cnt_reg_en;
wire [13:0] datain_w_cnt_st;
wire [13:0] datain_w_cnt_w;
wire [13:0] datain_w_cur;
wire datain_w_ori_reg_en;
wire [12:0] datain_width_cmp_w;
wire [13:0] datain_width_w;
wire [2:0] dataout_w_add;
wire [12:0] dataout_w_cnt_inc;
wire dataout_w_cnt_reg_en;
wire [12:0] dataout_w_cnt_w;
wire [12:0] dataout_w_init;
wire dataout_w_ori_reg_en;
wire [12:0] dataout_width_cmp_w;
wire [512 -1:0] dbg_csc_dat;
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: wire [8 -1:0] dbg_csc_dat_${i}; )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

wire [8 -1:0] dbg_csc_dat_0; 
wire [8 -1:0] dbg_csc_dat_1; 
wire [8 -1:0] dbg_csc_dat_2; 
wire [8 -1:0] dbg_csc_dat_3; 
wire [8 -1:0] dbg_csc_dat_4; 
wire [8 -1:0] dbg_csc_dat_5; 
wire [8 -1:0] dbg_csc_dat_6; 
wire [8 -1:0] dbg_csc_dat_7; 
wire [8 -1:0] dbg_csc_dat_8; 
wire [8 -1:0] dbg_csc_dat_9; 
wire [8 -1:0] dbg_csc_dat_10; 
wire [8 -1:0] dbg_csc_dat_11; 
wire [8 -1:0] dbg_csc_dat_12; 
wire [8 -1:0] dbg_csc_dat_13; 
wire [8 -1:0] dbg_csc_dat_14; 
wire [8 -1:0] dbg_csc_dat_15; 
wire [8 -1:0] dbg_csc_dat_16; 
wire [8 -1:0] dbg_csc_dat_17; 
wire [8 -1:0] dbg_csc_dat_18; 
wire [8 -1:0] dbg_csc_dat_19; 
wire [8 -1:0] dbg_csc_dat_20; 
wire [8 -1:0] dbg_csc_dat_21; 
wire [8 -1:0] dbg_csc_dat_22; 
wire [8 -1:0] dbg_csc_dat_23; 
wire [8 -1:0] dbg_csc_dat_24; 
wire [8 -1:0] dbg_csc_dat_25; 
wire [8 -1:0] dbg_csc_dat_26; 
wire [8 -1:0] dbg_csc_dat_27; 
wire [8 -1:0] dbg_csc_dat_28; 
wire [8 -1:0] dbg_csc_dat_29; 
wire [8 -1:0] dbg_csc_dat_30; 
wire [8 -1:0] dbg_csc_dat_31; 
wire [8 -1:0] dbg_csc_dat_32; 
wire [8 -1:0] dbg_csc_dat_33; 
wire [8 -1:0] dbg_csc_dat_34; 
wire [8 -1:0] dbg_csc_dat_35; 
wire [8 -1:0] dbg_csc_dat_36; 
wire [8 -1:0] dbg_csc_dat_37; 
wire [8 -1:0] dbg_csc_dat_38; 
wire [8 -1:0] dbg_csc_dat_39; 
wire [8 -1:0] dbg_csc_dat_40; 
wire [8 -1:0] dbg_csc_dat_41; 
wire [8 -1:0] dbg_csc_dat_42; 
wire [8 -1:0] dbg_csc_dat_43; 
wire [8 -1:0] dbg_csc_dat_44; 
wire [8 -1:0] dbg_csc_dat_45; 
wire [8 -1:0] dbg_csc_dat_46; 
wire [8 -1:0] dbg_csc_dat_47; 
wire [8 -1:0] dbg_csc_dat_48; 
wire [8 -1:0] dbg_csc_dat_49; 
wire [8 -1:0] dbg_csc_dat_50; 
wire [8 -1:0] dbg_csc_dat_51; 
wire [8 -1:0] dbg_csc_dat_52; 
wire [8 -1:0] dbg_csc_dat_53; 
wire [8 -1:0] dbg_csc_dat_54; 
wire [8 -1:0] dbg_csc_dat_55; 
wire [8 -1:0] dbg_csc_dat_56; 
wire [8 -1:0] dbg_csc_dat_57; 
wire [8 -1:0] dbg_csc_dat_58; 
wire [8 -1:0] dbg_csc_dat_59; 
wire [8 -1:0] dbg_csc_dat_60; 
wire [8 -1:0] dbg_csc_dat_61; 
wire [8 -1:0] dbg_csc_dat_62; 
wire [8 -1:0] dbg_csc_dat_63; 
//| eperl: generated_end (DO NOT EDIT ABOVE)
wire dl_block_end;
wire dl_channel_end;
wire [6:0] dl_channel_size;
wire [1:0] dl_cur_sub_h;
wire dl_dat_release;
wire dl_group_end;
wire [4:0] dl_h_offset;
wire [9:0] dl_h_offset_ext;
wire [30:0] dl_in_pd;
wire [30:0] dl_in_pd_d0;
wire dl_in_pvld;
wire dl_in_pvld_d0;
wire dl_layer_end;
wire [30:0] dl_pd;
wire [30:0] dl_pd_d0;
wire dl_pvld;
wire dl_pvld_d0;
wire [6:0] dl_stripe_length;
wire [4:0] dl_w_offset;
wire [9:0] dl_w_offset_ext;
wire [15 -1:0] entries_batch_w;
wire [15 -1:0] entries_single_w;
wire [15 -1:0] entries_w;
wire [13 -1:0] h_bias_0_stride_w;
wire [13 -1:0] h_bias_0_w;
wire [13 -1:0] h_bias_1_stride_w;
wire [13 -1:0] h_bias_1_w;
wire [13 -1:0] h_bias_2_w;
wire [13 -1:0] h_bias_3_w;
wire [13 -1:0] h_bias_d1;
wire [1:0] h_bias_reg_en;
wire [13:0] h_offset_slice_w;
wire is_batch_end;
wire is_conv;
wire is_dat_entry_end_wrap;
wire is_dat_entry_st_wrap;
wire is_dat_req_addr_wrap;
wire is_img;
wire is_last_channel;
wire is_pixel;
wire is_running_first;
wire is_sg_done;
wire is_sg_idle;
wire is_sg_running;
wire is_stripe_end;
wire is_stripe_equal;
wire is_sub_h_end;
wire is_w_end;
wire is_w_end_ahead;
wire is_winograd;
wire layer_st;
wire mon_batch_cnt_w;
wire mon_c_bias_w;
wire mon_dat_entry_avl_w;
wire mon_dat_entry_end_inc_wrap;
wire mon_dat_entry_st_inc_wrap;
wire [3:0] mon_dat_out_pra_vld;
wire [1:0] mon_dat_req_addr_wrap;
wire [512 -1:0] mon_dat_rsp_l0_sft;
wire [512 -1:0] mon_dat_rsp_l1_sft;
wire [512 -1:0] mon_dat_rsp_l2_sft;
wire [512 -1:0] mon_dat_rsp_l3_sft;
wire [3:0] mon_dat_rsp_pra_rdy;
wire mon_dat_slice_avl_w;
wire mon_data_bank_w;
wire mon_datain_c_cnt_inc;
wire mon_datain_h_cnt_inc;
wire mon_datain_h_cur;
wire mon_datain_w_cnt_inc;
wire mon_datain_w_cur;
wire mon_dataout_w_cnt_inc;
wire [5:0] mon_entries_batch_w;
wire mon_entries_single_w;
wire mon_entries_w;
wire [5:0] mon_h_bias_0_stride_w;
wire [13 -1:0] mon_h_bias_0_w;
wire [12:0] mon_h_bias_1_stride_w;
wire [4:0] mon_h_bias_1_w;
wire [4:0] mon_h_bias_2_w;
wire [1:0] mon_h_bias_3_w;
wire mon_h_bias_d1;
wire mon_pixel_w_cnt_w;
wire [1:0] mon_pixel_x_init_w;
wire mon_rls_slices_w;
wire mon_rsp_sft_cnt_l0_w;
wire mon_rsp_sft_cnt_l1_w;
wire mon_rsp_sft_cnt_l2_w;
wire mon_rsp_sft_cnt_l3_w;
wire [13:0] mon_slice_entries_w;
wire [1:0] mon_slice_left_w;
wire mon_stripe_cnt_inc;
wire [2:0] mon_sub_h_total_w;
wire pixel_ch_ori_reg_en;
wire [11:0] pixel_ch_stride_w;
wire pixel_force_clr;
wire pixel_force_fetch;
wire pixel_w_cnt_reg_en;
wire [15:0] pixel_w_cnt_w;
wire [14:0] pixel_w_cur;
wire pixel_w_ori_reg_en;
wire [7:0] pixel_x_add_w;
wire [6:0] pixel_x_byte_stride_w;
wire [6:0] pixel_x_cnt_add;
wire [6:0] pixel_x_init_offset_w;
wire [5:0] pixel_x_init_w;
wire [5:0] pixel_x_stride_w;
wire [1:0] pra_precision_0;
wire [1:0] pra_precision_1;
wire [1:0] pra_precision_2;
wire [1:0] pra_precision_3;
wire [1:0] pra_truncate_0;
wire [1:0] pra_truncate_1;
wire [1:0] pra_truncate_2;
wire [1:0] pra_truncate_3;
wire [1:0] pra_truncate_w;
wire reuse_rls;
wire [13:0] rls_slices_w;
wire rsp_sft_cnt_l0_en;
wire [7:0] rsp_sft_cnt_l0_inc;
wire rsp_sft_cnt_l0_ori_en;
wire [7:0] rsp_sft_cnt_l0_sub;
wire [7:0] rsp_sft_cnt_l0_w;
wire rsp_sft_cnt_l1_en;
wire [7:0] rsp_sft_cnt_l1_inc;
wire rsp_sft_cnt_l1_ori_en;
wire [7:0] rsp_sft_cnt_l1_sub;
wire [7:0] rsp_sft_cnt_l1_w;
wire rsp_sft_cnt_l2_en;
wire [7:0] rsp_sft_cnt_l2_inc;
wire rsp_sft_cnt_l2_ori_en;
wire [7:0] rsp_sft_cnt_l2_sub;
wire [7:0] rsp_sft_cnt_l2_w;
wire rsp_sft_cnt_l3_en;
wire [7:0] rsp_sft_cnt_l3_inc;
wire rsp_sft_cnt_l3_ori_en;
wire [7:0] rsp_sft_cnt_l3_sub;
wire [7:0] rsp_sft_cnt_l3_w;
wire rsp_sft_l1_sel_1;
wire rsp_sft_l1_sel_2;
wire rsp_sft_l1_sel_3;
wire rsp_sft_l2_sel_1;
wire rsp_sft_l2_sel_2;
wire rsp_sft_l2_sel_3;
wire rsp_sft_l3_sel_1;
wire rsp_sft_l3_sel_2;
wire rsp_sft_l3_sel_3;
wire sc2buf_dat_rd_en_w;
wire [15 -1:0] sc2cdma_dat_entries_w;
wire [13:0] sc2cdma_dat_slices_w;
wire [8:0] sc2mac_dat_pd_w;
wire slcg_wg_en_w;
wire [15 -1:0] slice_entries_w;
wire [13:0] slice_left_w;
wire [13:0] slices_oprand;
wire [6:0] stripe_cnt_inc;
wire stripe_cnt_reg_en;
wire [6:0] stripe_cnt_w;
wire [2:0] sub_h_cmp_w;
wire [2:0] sub_h_cnt_inc;
wire sub_h_cnt_reg_en;
wire [1:0] sub_h_cnt_w;
wire [2:0] sub_h_total_w;
wire sub_rls;
wire [14:0] w_bias_int8;
wire w_bias_reg_en;
wire [13:0] w_bias_w;
wire [5:0] x_dilate_w;
wire [5:0] y_dilate_w;
/////////////////////////////////////////////////////////////////////////////////////////////
// Pipeline of Weight loader, for both compressed weight and uncompressed weight
//
// input_package
// |
// data request
// |
// conv_buffer
// |
// feature data---> data relase
// | |
// REG PRA
// | |
// REGISTER
// |
// MAC
//
/////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////
///// status from sequence generator                     /////
//////////////////////////////////////////////////////////////
assign is_sg_idle = (sc_state == 0 );
assign is_sg_running = (sc_state == 2 );
assign is_sg_done = (sc_state == 3 );
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"is_sg_running\" -q is_sg_running_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       is_sg_running_d1 <= 1'b0;
   end else begin
       is_sg_running_d1 <= is_sg_running;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// input signals from registers                       /////
//////////////////////////////////////////////////////////////
assign layer_st = reg2dp_op_en & is_sg_idle;
assign is_pixel = (reg2dp_datain_format == 1'h1 );
assign is_winograd = 1'b0;
assign is_conv = (reg2dp_conv_mode == 1'h0 );
assign is_img = is_conv & is_pixel;
assign {mon_data_bank_w, data_bank_w} = reg2dp_data_bank + 1'b1;
assign data_batch_w = 6'b1;
assign batch_cmp_w = 5'b0;
//assign is_int8 = (reg2dp_proc_precision == 2'h0 );
//assign is_fp16 = (reg2dp_proc_precision == 2'h2 );
assign datain_width_w = is_winograd ? ({2'b0, reg2dp_datain_width_ext[12:2]} + 1'b1) : reg2dp_datain_width_ext + 1'b1;
assign datain_width_cmp_w = reg2dp_datain_width_ext;
assign datain_height_cmp_w = reg2dp_datain_height_ext;
assign datain_channel_cmp_w = is_winograd ? reg2dp_weight_channel_ext[12:2] : {{6 -2{1'b0}}, reg2dp_weight_channel_ext[12:6]};
//y_ex=0,sub_h_total=1;y_ex=1,sub_h_total=2; y_ext=2,sub_h_total=4; non_image, sub_h_total=1;
//sub_h_total means how many h lines are used in post-extention
assign {sub_h_total_w, mon_sub_h_total_w} = is_img ? (6'h9 << reg2dp_y_extension) : 6'h8;
assign sub_h_cmp_w = is_img ? sub_h_total_w : is_winograd ? 3'h2 : 3'h1;
assign dataout_w_init[12:0] = sub_h_cmp_w - 1'b1;
assign conv_x_stride_w = (is_winograd) ? 4'b1 : reg2dp_conv_x_stride_ext + 1'b1;
assign pixel_x_stride_w = (reg2dp_datain_channel_ext[1:0] == 2'h3) ? {conv_x_stride_w, 2'b0} : //*4, after pre_extension
                          (reg2dp_datain_channel_ext[1:0] == 2'h2) ? ({conv_x_stride_w, 1'b0} + conv_x_stride_w) : //*3
                          {2'b0, conv_x_stride_w}; //*1
//: my $kk=6;
//: if ($kk=6) {
//: print qq (
//: assign {mon_pixel_x_init_w,pixel_x_init_w} = (reg2dp_y_extension == 2'h2) ? ({pixel_x_stride_w, 1'b0} + pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]) :
//: (reg2dp_y_extension == 2'h1) ? (pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]):
//: (reg2dp_weight_channel_ext >= 7'h40) ? {6{1'b1}}: //cut by atomC
//: {reg2dp_weight_channel_ext[6 -1:0]};
//: )
//: }
//: else {
//: print qq(
//: assign {mon_pixel_x_init_w,pixel_x_init_w} = (reg2dp_y_extension == 2'h2) ? ({pixel_x_stride_w, 1'b0} + pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]) :
//: (reg2dp_y_extension == 2'h1) ? (pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]):
//: (reg2dp_weight_channel_ext >= 7'h40) ? {6{1'b1}}: //cut by atomC
//: {{6-6{1'b0}},reg2dp_weight_channel_ext[6 -1:0]};
//: )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

assign {mon_pixel_x_init_w,pixel_x_init_w} = (reg2dp_y_extension == 2'h2) ? ({pixel_x_stride_w, 1'b0} + pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]) :
(reg2dp_y_extension == 2'h1) ? (pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]):
(reg2dp_weight_channel_ext >= 7'h40) ? {6{1'b1}}: //cut by atomC
{reg2dp_weight_channel_ext[6 -1:0]};

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign pixel_x_init_offset_w = (reg2dp_weight_channel_ext[6 -1:0] + 1'b1);
assign pixel_x_add_w = (reg2dp_y_extension == 2'h2) ? {pixel_x_stride_w, 2'b0} : //*4, after post_extension
                       (reg2dp_y_extension == 2'h1) ? {1'b0, pixel_x_stride_w, 1'b0} : //*2
                       {2'b0, pixel_x_stride_w};
assign pixel_x_byte_stride_w = {1'b0, pixel_x_stride_w};
//: my $kk=5;
//: if($kk=5) {
//: print qq(
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_1
//: assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_2
//: assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_4
//: assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +2{1'b0}}}; //stick to 4*atomK  no matter which config.  
//: `endif
//: )
//: }
//: else {
//: print qq(
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_1
//: assign pixel_ch_stride_w = {{5-5{1'b0}},pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_2
//: assign pixel_ch_stride_w = {{5-5{1'b0}},pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_4
//: assign pixel_ch_stride_w = {{5-5{1'b0}},pixel_x_stride_w, {5 +2{1'b0}}}; //stick to 4*atomK  no matter which config.  
//: `endif
//: )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  


//| eperl: generated_end (DO NOT EDIT ABOVE)
assign conv_y_stride_w = (is_winograd) ? 4'b1 : reg2dp_conv_y_stride_ext + 1'b1;
assign x_dilate_w = (is_winograd | is_img) ? 6'b1 : reg2dp_x_dilation_ext + 1'b1;
assign y_dilate_w = (is_winograd | is_img) ? 6'b1 : reg2dp_y_dilation_ext + 1'b1;
//reg2dp_entries means entry per slice
assign {mon_entries_single_w,entries_single_w} = (reg2dp_entries + 1'b1);
assign {mon_entries_batch_w,entries_batch_w} = entries_single_w * data_batch_w;
assign {mon_entries_w,entries_w} = (is_winograd) ? ({reg2dp_entries[12:0], 2'b0} + 3'h4) : entries_single_w;
assign h_offset_slice_w[11:0] = data_batch_w * y_dilate_w;
assign h_offset_slice_w[13:12] = 2'b0;
assign {mon_h_bias_0_stride_w,h_bias_0_stride_w} = entries * data_batch;
assign {mon_h_bias_1_stride_w,h_bias_1_stride_w} = entries * h_offset_slice;
assign {mon_rls_slices_w,rls_slices_w} = reg2dp_rls_slices + 1'b1;
assign {mon_slice_left_w,slice_left_w} = reg2dp_skip_data_rls ? (reg2dp_datain_height_ext + 1'b1) : reg2dp_datain_height_ext - reg2dp_rls_slices;
assign slices_oprand = layer_st_d1 ? rls_slices : slice_left;
assign {mon_slice_entries_w,slice_entries_w} = entries_batch * slices_oprand;
assign dataout_width_cmp_w = reg2dp_dataout_width;
assign pra_truncate_w = (reg2dp_pra_truncate == 2'h3) ? 2'h2 : reg2dp_pra_truncate;
//: my $kk=15;
//: my $jj=13;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"layer_st\" -q layer_st_d1");
//: &eperl::flop("-nodeclare   -rval \"{22{1'b0}}\"  -en \"layer_st\" -d \"{22{is_winograd}}\" -q is_winograd_d1");
//: &eperl::flop("-nodeclare   -rval \"{34{1'b0}}\"  -en \"layer_st\" -d \"{34{is_img}}\" -q is_img_d1");
//: &eperl::flop("-nodeclare   -rval \"{5{1'b0}}\"  -en \"layer_st\" -d \"data_bank_w\" -q data_bank");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"datain_width_w\" -q datain_width");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"layer_st\" -d \"datain_width_cmp_w\" -q datain_width_cmp");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"layer_st\" -d \"datain_height_cmp_w\" -q datain_height_cmp");
//: &eperl::flop("-nodeclare   -rval \"{11{1'b0}}\"  -en \"layer_st\" -d \"datain_channel_cmp_w\" -q datain_channel_cmp");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g0");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g1");
//: &eperl::flop("-nodeclare   -rval \"2'h1\"  -en \"layer_st\" -d \"sub_h_total_w[2:1]\" -q sub_h_total_g2");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g3");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g4");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g5");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g6");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g7");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g8");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g9");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g10");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g11");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_cmp_w\" -q sub_h_cmp_g0");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_cmp_w\" -q sub_h_cmp_g1");
//: &eperl::flop("-nodeclare   -rval \"{4{1'b0}}\"  -en \"layer_st\" -d \"conv_x_stride_w\" -q conv_x_stride");
//: &eperl::flop("-nodeclare   -rval \"{4{1'b0}}\"  -en \"layer_st\" -d \"conv_y_stride_w\" -q conv_y_stride");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"layer_st\" -d \"pixel_x_stride_w[0]\" -q pixel_x_stride_odd");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"data_batch_w\" -q data_batch");
//: &eperl::flop("-nodeclare   -rval \"{5{1'b0}}\"  -en \"layer_st\" -d \"batch_cmp_w\" -q batch_cmp");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_init_w\" -q pixel_x_init");
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_init_offset_w\" -q pixel_x_init_offset");
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_add_w[6:0]\" -q pixel_x_add");
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_byte_stride_w\" -q pixel_x_byte_stride");
//: &eperl::flop("-nodeclare   -rval \"{12{1'b0}}\"  -en \"layer_st\" -d \"pixel_ch_stride_w\" -q pixel_ch_stride");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"x_dilate_w\" -q x_dilate");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"y_dilate_w\" -q y_dilate");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"layer_st\" -d \"reg2dp_pad_value\" -q pad_value");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st\" -d \"entries_w\" -q entries");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st\" -d \"entries_batch_w\" -q entries_batch");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st\" -d \"{1'h0,reg2dp_entries}\" -q entries_cmp");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"h_offset_slice_w\" -q h_offset_slice");
//: &eperl::flop("-nodeclare   -rval \"{12{1'b0}}\"  -en \"layer_st_d1\" -d \"h_bias_0_stride_w\" -q h_bias_0_stride");
//: &eperl::flop("-nodeclare   -rval \"{12{1'b0}}\"  -en \"layer_st_d1\" -d \"h_bias_1_stride_w\" -q h_bias_1_stride");
//: &eperl::flop("-nodeclare   -rval \"{${jj}{1'b0}}\"  -en \"layer_st_d1\" -d \"entries[${jj}-1:0]\" -q h_bias_2_stride");
//: &eperl::flop("-nodeclare   -rval \"{${jj}{1'b0}}\"  -en \"layer_st_d1\" -d \"entries[${jj}-1:0]\" -q h_bias_3_stride");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"rls_slices_w\" -q rls_slices");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st_d1\" -d \"slice_entries_w\" -q rls_entries");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"slice_left_w[13:0]\" -q slice_left");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"is_sg_done\" -d \"slice_left\" -q last_slices");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"is_sg_done\" -d \"slice_entries_w\" -q last_entries");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"layer_st\" -d \"dataout_width_cmp_w\" -q dataout_width_cmp");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"layer_st\" -d \"{4{pra_truncate_w}}\" -q pra_truncate");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"layer_st\" -d \"{4{reg2dp_proc_precision}}\" -q pra_precision");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       layer_st_d1 <= 1'b0;
   end else begin
       layer_st_d1 <= layer_st;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       is_winograd_d1 <= {22{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           is_winograd_d1 <= {22{is_winograd}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           is_winograd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       is_img_d1 <= {34{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           is_img_d1 <= {34{is_img}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           is_img_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       data_bank <= {5{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           data_bank <= data_bank_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           data_bank <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_width <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_width <= datain_width_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_width <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_width_cmp <= {13{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_width_cmp <= datain_width_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_width_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_height_cmp <= {13{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_height_cmp <= datain_height_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_height_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_channel_cmp <= {11{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_channel_cmp <= datain_channel_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_channel_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g0 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g0 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g0 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g1 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g1 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g2 <= 2'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g2 <= sub_h_total_w[2:1];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g3 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g3 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g4 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g4 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g4 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g5 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g5 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g5 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g6 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g6 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g6 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g7 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g7 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g7 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g8 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g8 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g8 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g9 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g9 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g9 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g10 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g10 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g10 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g11 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g11 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g11 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_cmp_g0 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_cmp_g0 <= sub_h_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_cmp_g0 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_cmp_g1 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_cmp_g1 <= sub_h_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_cmp_g1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       conv_x_stride <= {4{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           conv_x_stride <= conv_x_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           conv_x_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       conv_y_stride <= {4{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           conv_y_stride <= conv_y_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           conv_y_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_stride_odd <= 1'b0;
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_stride_odd <= pixel_x_stride_w[0];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_stride_odd <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       data_batch <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           data_batch <= data_batch_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           data_batch <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       batch_cmp <= {5{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           batch_cmp <= batch_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           batch_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_init <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_init <= pixel_x_init_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_init <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_init_offset <= {7{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_init_offset <= pixel_x_init_offset_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_init_offset <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_add <= {7{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_add <= pixel_x_add_w[6:0];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_add <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_byte_stride <= {7{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_byte_stride <= pixel_x_byte_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_byte_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_ch_stride <= {12{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_ch_stride <= pixel_ch_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_ch_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       x_dilate <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           x_dilate <= x_dilate_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           x_dilate <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       y_dilate <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           y_dilate <= y_dilate_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           y_dilate <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pad_value <= {16{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pad_value <= reg2dp_pad_value;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pad_value <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       entries <= {15{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           entries <= entries_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           entries <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       entries_batch <= {15{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           entries_batch <= entries_batch_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           entries_batch <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       entries_cmp <= {15{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           entries_cmp <= {1'h0,reg2dp_entries};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           entries_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_offset_slice <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           h_offset_slice <= h_offset_slice_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           h_offset_slice <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_0_stride <= {12{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_0_stride <= h_bias_0_stride_w;
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_0_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_1_stride <= {12{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_1_stride <= h_bias_1_stride_w;
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_1_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_2_stride <= {13{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_2_stride <= entries[13-1:0];
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_2_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_3_stride <= {13{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_3_stride <= entries[13-1:0];
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_3_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rls_slices <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           rls_slices <= rls_slices_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           rls_slices <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rls_entries <= {15{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           rls_entries <= slice_entries_w;
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           rls_entries <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slice_left <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           slice_left <= slice_left_w[13:0];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           slice_left <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       last_slices <= {14{1'b0}};
   end else begin
       if ((is_sg_done) == 1'b1) begin
           last_slices <= slice_left;
       // VCS coverage off
       end else if ((is_sg_done) == 1'b0) begin
       end else begin
           last_slices <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       last_entries <= {15{1'b0}};
   end else begin
       if ((is_sg_done) == 1'b1) begin
           last_entries <= slice_entries_w;
       // VCS coverage off
       end else if ((is_sg_done) == 1'b0) begin
       end else begin
           last_entries <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dataout_width_cmp <= {13{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           dataout_width_cmp <= dataout_width_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           dataout_width_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pra_truncate <= {8{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pra_truncate <= {4{pra_truncate_w}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pra_truncate <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pra_precision <= {8{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pra_precision <= {4{reg2dp_proc_precision}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pra_precision <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////////////////////////////////////////////////////
// SLCG control signal //
////////////////////////////////////////////////////////////////////////
assign slcg_wg_en_w = reg2dp_op_en & is_winograd;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"slcg_wg_en_w\" -q slcg_wg_en_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"slcg_wg_en_d1\" -q slcg_wg_en_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"slcg_wg_en_d2\" -q slcg_wg_en_d3");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slcg_wg_en_d1 <= 1'b0;
   end else begin
       slcg_wg_en_d1 <= slcg_wg_en_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slcg_wg_en_d2 <= 1'b0;
   end else begin
       slcg_wg_en_d2 <= slcg_wg_en_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slcg_wg_en_d3 <= 1'b0;
   end else begin
       slcg_wg_en_d3 <= slcg_wg_en_d2;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign slcg_wg_en = slcg_wg_en_d3;
//////////////////////////////////////////////////////////////
///// cbuf status management                             /////
//////////////////////////////////////////////////////////////
//================ Non-SLCG clock domain ================//
assign cbuf_reset = sc2cdma_dat_pending_req;
assign is_running_first = is_sg_running & ~is_sg_running_d1;
//////////////////////////////////// calculate how many avaliable dat slices in cbuf////////////////////////////////////
assign dat_slice_avl_add = cdma2sc_dat_updt ? cdma2sc_dat_slices : 14'b0;
assign dat_slice_avl_sub = dat_rls ? sc2cdma_dat_slices_w : 14'b0;
assign {mon_dat_slice_avl_w, dat_slice_avl_w} = (cbuf_reset) ? 14'b0 : dat_slice_avl + dat_slice_avl_add - dat_slice_avl_sub;
//////////////////////////////////// calculate how many avaliable dat entries in cbuf////////////////////////////////////
assign dat_entry_avl_add = cdma2sc_dat_updt ? cdma2sc_dat_entries :{15{1'b0}};
assign dat_entry_avl_sub = dat_rls ? sc2cdma_dat_entries_w : {15{1'b0}};
assign {mon_dat_entry_avl_w,dat_entry_avl_w} = (cbuf_reset) ? {15{1'b0}} : dat_entry_avl + dat_entry_avl_add - dat_entry_avl_sub;
//////////////////////////////////// calculate avilable data entries start offset in cbuf banks ////////////////////////////////////
// data_bank is the highest bank for storing data
assign {mon_dat_entry_st_inc,dat_entry_st_inc} = dat_entry_st + dat_entry_avl_sub;
assign {mon_dat_entry_st_inc_wrap, dat_entry_st_inc_wrap} = dat_entry_st_inc - {data_bank, {9{1'b0}} };
assign is_dat_entry_st_wrap = (dat_entry_st_inc >= {1'b0, data_bank, {9{1'b0}} });
assign dat_entry_st_w = (cbuf_reset) ? {15{1'b0}} : is_dat_entry_st_wrap ? dat_entry_st_inc_wrap : dat_entry_st_inc[15 -1:0];
//////////////////////////////////// calculate avilable data entries end offset in cbuf banks////////////////////////////////////
assign {mon_dat_entry_end_inc,dat_entry_end_inc} = dat_entry_end + dat_entry_avl_add;
assign {mon_dat_entry_end_inc_wrap,dat_entry_end_inc_wrap} = dat_entry_end_inc - {data_bank, {9{1'b0}} };
assign is_dat_entry_end_wrap = (dat_entry_end_inc >= {1'b0, data_bank, {9{1'b0}} });
assign dat_entry_end_w = (cbuf_reset) ? {15{1'b0}} : is_dat_entry_end_wrap ? dat_entry_end_inc_wrap : dat_entry_end_inc[15 -1:0];
//////////////////////////////////// registers and assertions ////////////////////////////////////
//: my $kk= 15;
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{14{1'b0}}\"  -en \"cdma2sc_dat_updt | dat_rls | cbuf_reset\" -d \"dat_slice_avl_w\" -q dat_slice_avl");
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{${kk}{1'b0}}\"  -en \"cdma2sc_dat_updt | dat_rls | cbuf_reset\" -d \"dat_entry_avl_w\" -q dat_entry_avl");
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{${kk}{1'b0}}\"  -en \"cbuf_reset | dat_rls\" -d \"dat_entry_st_w\" -q dat_entry_st");
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{${kk}{1'b0}}\"  -en \"cbuf_reset | cdma2sc_dat_updt\" -d \"dat_entry_end_w\" -q dat_entry_end");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_ng_clk or negedge nvdla_core_rstn) begin
   if (!nvdla_core_rstn) begin
       dat_slice_avl <= {14{1'b0}};
   end else begin
       if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b1) begin
           dat_slice_avl <= dat_slice_avl_w;
       // VCS coverage off
       end else if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b0) begin
       end else begin
           dat_slice_avl <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_ng_clk or negedge nvdla_core_rstn) begin
   if (!nvdla_core_rstn) begin
       dat_entry_avl <= {15{1'b0}};
   end else begin
       if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b1) begin
           dat_entry_avl <= dat_entry_avl_w;
       // VCS coverage off
       end else if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b0) begin
       end else begin
           dat_entry_avl <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_ng_clk or negedge nvdla_core_rstn) begin
   if (!nvdla_core_rstn) begin
       dat_entry_st <= {15{1'b0}};
   end else begin
       if ((cbuf_reset | dat_rls) == 1'b1) begin
           dat_entry_st <= dat_entry_st_w;
       // VCS coverage off
       end else if ((cbuf_reset | dat_rls) == 1'b0) begin
       end else begin
           dat_entry_st <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_ng_clk or negedge nvdla_core_rstn) begin
   if (!nvdla_core_rstn) begin
       dat_entry_end <= {15{1'b0}};
   end else begin
       if ((cbuf_reset | cdma2sc_dat_updt) == 1'b1) begin
           dat_entry_end <= dat_entry_end_w;
       // VCS coverage off
       end else if ((cbuf_reset | cdma2sc_dat_updt) == 1'b0) begin
       end else begin
           dat_entry_end <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//================ Non-SLCG clock domain end ================//
//////////////////////////////////////////////////////////////
///// cbuf status update                                 /////
//////////////////////////////////////////////////////////////
assign sub_rls = (dat_rsp_pvld & dat_rsp_rls);
assign reuse_rls = sg2dl_reuse_rls;
assign dat_rls = (reuse_rls & (|last_slices)) | (sub_rls & (|rls_slices));
assign sc2cdma_dat_slices_w = sub_rls ? rls_slices : last_slices;
assign sc2cdma_dat_entries_w = sub_rls ? rls_entries : last_entries;
//: my $kk=15;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_rls\" -q sc2cdma_dat_updt");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"dat_rls\" -d \"sc2cdma_dat_slices_w[13:0]\" -q sc2cdma_dat_slices");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dat_rls\" -d \"sc2cdma_dat_entries_w\" -q sc2cdma_dat_entries");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2cdma_dat_updt <= 1'b0;
   end else begin
       sc2cdma_dat_updt <= dat_rls;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2cdma_dat_slices <= {14{1'b0}};
   end else begin
       if ((dat_rls) == 1'b1) begin
           sc2cdma_dat_slices <= sc2cdma_dat_slices_w[13:0];
       // VCS coverage off
       end else if ((dat_rls) == 1'b0) begin
       end else begin
           sc2cdma_dat_slices <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2cdma_dat_entries <= {15{1'b0}};
   end else begin
       if ((dat_rls) == 1'b1) begin
           sc2cdma_dat_entries <= sc2cdma_dat_entries_w;
       // VCS coverage off
       end else if ((dat_rls) == 1'b0) begin
       end else begin
           sc2cdma_dat_entries <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// input sg2dl package                                 /////
//////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////
///// generate data read sequence                        /////
//////////////////////////////////////////////////////////////
//: my $total_depth = 0 + 5;
//: my $wg_depth = 0;
//:
//: print "assign dl_in_pvld_d0 = sg2dl_pvld;\n";
//: print "assign dl_in_pd_d0 = sg2dl_pd;\n\n";
//:
//: for(my $i = 0; $i < $total_depth; $i ++) {
//: my $j = $i + 1;
//: &eperl::flop("-wid 1    -rval \"1'b0\"                                 -d \"dl_in_pvld_d${i}\" -q dl_in_pvld_d${j}");
//: &eperl::flop("-wid 31   -rval \"{31{1'b0}}\"  -en \"dl_in_pvld_d${i}\" -d \"dl_in_pd_d${i}\"   -q dl_in_pd_d${j}");
//: }
//:
//: my $d0 = $total_depth;
//: my $d1 = $wg_depth;
//:
//: print "assign dl_in_pvld = (is_winograd_d1[0]) ? dl_in_pvld_d${d1} : dl_in_pvld_d${d0};\n";
//: print "assign dl_in_pd = (is_winograd_d1[1]) ? dl_in_pd_d${d1} : dl_in_pd_d${d0};\n\n";
//: my $pipe_depth = 4;
//: my $i;
//: my $j;
//: print "assign dl_pvld_d0 = dl_in_pvld;\n";
//: print "assign dl_pd_d0 = dl_in_pd;\n\n";
//: for($i = 0; $i < $pipe_depth; $i ++) {
//: $j = $i + 1;
//: &eperl::flop("-nodeclare -rval \"1'b0\"                              -d \"dl_pvld_d${i}\"   -q dl_pvld_d${j}");
//: &eperl::flop("-nodeclare -rval \"{31{1'b0}}\"  -en \"dl_pvld_d${i}\" -d \"dl_pd_d${i}\"     -q dl_pd_d${j}");
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dl_in_pvld_d0 = sg2dl_pvld;
assign dl_in_pd_d0 = sg2dl_pd;

reg  dl_in_pvld_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d1 <= 1'b0;
   end else begin
       dl_in_pvld_d1 <= dl_in_pvld_d0;
   end
end
reg [30:0] dl_in_pd_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d1 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d0) == 1'b1) begin
           dl_in_pd_d1 <= dl_in_pd_d0;
       // VCS coverage off
       end else if ((dl_in_pvld_d0) == 1'b0) begin
       end else begin
           dl_in_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d2 <= 1'b0;
   end else begin
       dl_in_pvld_d2 <= dl_in_pvld_d1;
   end
end
reg [30:0] dl_in_pd_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d2 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d1) == 1'b1) begin
           dl_in_pd_d2 <= dl_in_pd_d1;
       // VCS coverage off
       end else if ((dl_in_pvld_d1) == 1'b0) begin
       end else begin
           dl_in_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d3 <= 1'b0;
   end else begin
       dl_in_pvld_d3 <= dl_in_pvld_d2;
   end
end
reg [30:0] dl_in_pd_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d3 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d2) == 1'b1) begin
           dl_in_pd_d3 <= dl_in_pd_d2;
       // VCS coverage off
       end else if ((dl_in_pvld_d2) == 1'b0) begin
       end else begin
           dl_in_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d4 <= 1'b0;
   end else begin
       dl_in_pvld_d4 <= dl_in_pvld_d3;
   end
end
reg [30:0] dl_in_pd_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d4 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d3) == 1'b1) begin
           dl_in_pd_d4 <= dl_in_pd_d3;
       // VCS coverage off
       end else if ((dl_in_pvld_d3) == 1'b0) begin
       end else begin
           dl_in_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d5 <= 1'b0;
   end else begin
       dl_in_pvld_d5 <= dl_in_pvld_d4;
   end
end
reg [30:0] dl_in_pd_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d5 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d4) == 1'b1) begin
           dl_in_pd_d5 <= dl_in_pd_d4;
       // VCS coverage off
       end else if ((dl_in_pvld_d4) == 1'b0) begin
       end else begin
           dl_in_pd_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
assign dl_in_pvld = (is_winograd_d1[0]) ? dl_in_pvld_d0 : dl_in_pvld_d5;
assign dl_in_pd = (is_winograd_d1[1]) ? dl_in_pd_d0 : dl_in_pd_d5;

assign dl_pvld_d0 = dl_in_pvld;
assign dl_pd_d0 = dl_in_pd;

always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d1 <= 1'b0;
   end else begin
       dl_pvld_d1 <= dl_pvld_d0;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d1 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d0) == 1'b1) begin
           dl_pd_d1 <= dl_pd_d0;
       // VCS coverage off
       end else if ((dl_pvld_d0) == 1'b0) begin
       end else begin
           dl_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d2 <= 1'b0;
   end else begin
       dl_pvld_d2 <= dl_pvld_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d2 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d1) == 1'b1) begin
           dl_pd_d2 <= dl_pd_d1;
       // VCS coverage off
       end else if ((dl_pvld_d1) == 1'b0) begin
       end else begin
           dl_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d3 <= 1'b0;
   end else begin
       dl_pvld_d3 <= dl_pvld_d2;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d3 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d2) == 1'b1) begin
           dl_pd_d3 <= dl_pd_d2;
       // VCS coverage off
       end else if ((dl_pvld_d2) == 1'b0) begin
       end else begin
           dl_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d4 <= 1'b0;
   end else begin
       dl_pvld_d4 <= dl_pvld_d3;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d4 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d3) == 1'b1) begin
           dl_pd_d4 <= dl_pd_d3;
       // VCS coverage off
       end else if ((dl_pvld_d3) == 1'b0) begin
       end else begin
           dl_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dl_pvld = (sub_h_total_g0[2] & dl_pvld_d1) |
                 (sub_h_total_g0[1] & dl_pvld_d3) |
                 (sub_h_total_g0[0] & dl_pvld_d4);
assign dl_pd = ({31 {sub_h_total_g1[2]}} & dl_pd_d1) |
               ({31 {sub_h_total_g1[1]}} & dl_pd_d3) |
               ({31 {sub_h_total_g1[0]}} & dl_pd_d4);
// PKT_UNPACK_WIRE( csc_dat_pkg , dl_ , dl_pd )
assign dl_w_offset[4:0] = dl_pd[4:0]; //this is weight offset
assign dl_h_offset[4:0] = dl_pd[9:5]; //weight offset
assign dl_channel_size[6:0] = dl_pd[16:10];
assign dl_stripe_length[6:0]= dl_pd[23:17];
assign dl_cur_sub_h[1:0] = dl_pd[25:24];
assign dl_block_end = dl_pd[26];
assign dl_channel_end = dl_pd[27];
assign dl_group_end = dl_pd[28];
assign dl_layer_end = dl_pd[29];
assign dl_dat_release = dl_pd[30];
////////////////////////// batch up counter //////////////////////////
assign {mon_batch_cnt_w,batch_cnt_w} = layer_st ? 6'b0 : is_batch_end ? 6'b0 : batch_cnt + 1'b1;
assign is_batch_end = (batch_cnt == batch_cmp);
//: &eperl::flop("-nodeclare   -rval \"{5{1'b0}}\"  -en \"layer_st | dat_exec_valid\" -d \"batch_cnt_w\" -q batch_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       batch_cnt <= {5{1'b0}};
   end else begin
       if ((layer_st | dat_exec_valid) == 1'b1) begin
           batch_cnt <= batch_cnt_w;
       // VCS coverage off
       end else if ((layer_st | dat_exec_valid) == 1'b0) begin
       end else begin
           batch_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// sub height up counter //////////////////////////
assign sub_h_cnt_inc = sub_h_cnt + 1'b1;
assign sub_h_cnt_w = (layer_st | is_sub_h_end) ? 2'b0 : sub_h_cnt_inc[1:0];
assign is_sub_h_end = (sub_h_cnt_inc == sub_h_cmp_g0);
assign sub_h_cnt_reg_en = layer_st | ((is_winograd_d1[2] | (|reg2dp_y_extension)) & dat_exec_valid);
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"sub_h_cnt_reg_en\" -d \"sub_h_cnt_w\" -q sub_h_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_cnt <= {2{1'b0}};
   end else begin
       if ((sub_h_cnt_reg_en) == 1'b1) begin
           sub_h_cnt <= sub_h_cnt_w;
       // VCS coverage off
       end else if ((sub_h_cnt_reg_en) == 1'b0) begin
       end else begin
           sub_h_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// stripe up counter //////////////////////////
assign {mon_stripe_cnt_inc,stripe_cnt_inc} = stripe_cnt + 1'b1;
assign stripe_cnt_w = layer_st ? 7'b0 :
                      (is_stripe_equal & ~is_sub_h_end) ? stripe_cnt :
                      is_stripe_end ? 7'b0 :
                      stripe_cnt_inc;
assign is_stripe_equal = is_batch_end & (stripe_cnt_inc == dl_stripe_length);
assign is_stripe_end = is_stripe_equal & is_sub_h_end;
assign stripe_cnt_reg_en = layer_st | (dat_exec_valid & is_batch_end);
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"stripe_cnt_reg_en\" -d \"stripe_cnt_w\" -q stripe_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       stripe_cnt <= {7{1'b0}};
   end else begin
       if ((stripe_cnt_reg_en) == 1'b1) begin
           stripe_cnt <= stripe_cnt_w;
       // VCS coverage off
       end else if ((stripe_cnt_reg_en) == 1'b0) begin
       end else begin
           stripe_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// pipe valid generator //////////////////////////
assign dat_pipe_local_valid_w = (dat_pipe_valid & is_stripe_equal) ? 1'b0 : dl_pvld ? 1'b1 : dat_pipe_local_valid;
assign dat_pipe_valid = dl_pvld | dat_pipe_local_valid;
assign dat_exec_valid = dl_pvld ? 1'b1 : (~(|stripe_cnt) & ~(|sub_h_cnt) & ~(|batch_cnt)) ? 1'b0 : dat_exec_valid_d1;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_pipe_local_valid_w\" -q dat_pipe_local_valid");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_pipe_valid\" -q dat_pipe_valid_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_exec_valid\" -q dat_exec_valid_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_pipe_local_valid <= 1'b0;
   end else begin
       dat_pipe_local_valid <= dat_pipe_local_valid_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_pipe_valid_d1 <= 1'b0;
   end else begin
       dat_pipe_valid_d1 <= dat_pipe_valid;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_exec_valid_d1 <= 1'b0;
   end else begin
       dat_exec_valid_d1 <= dat_exec_valid;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// request bytes //////////////////////////
assign dat_req_bytes = {1'b0, dl_channel_size};
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"dat_exec_valid\" -d \"dat_req_bytes\" -q dat_req_bytes_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_bytes_d1 <= {8{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_bytes_d1 <= dat_req_bytes;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_bytes_d1 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// output width coordinate counter //////////////////////////
// sub_h T, output will compute sub_h point in w direction
assign dataout_w_add = sub_h_cmp_g1;
assign {mon_dataout_w_cnt_inc,dataout_w_cnt_inc} = dataout_w_cnt + dataout_w_add;
assign is_w_end = is_batch_end & is_sub_h_end & (dataout_w_cnt >= dataout_width_cmp);
assign is_w_end_ahead = is_batch_end & (dataout_w_cnt >= dataout_width_cmp);
assign dataout_w_cnt_w = layer_st ? dataout_w_init :
                         (is_stripe_end & ~dl_channel_end) ? dataout_w_ori :
                         is_w_end ? dataout_w_init :
                         dataout_w_cnt_inc;
assign dataout_w_cnt_reg_en = layer_st | (dat_exec_valid & is_batch_end & is_sub_h_end);
assign dataout_w_ori_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_channel_end);
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"dataout_w_cnt_reg_en\" -d \"dataout_w_cnt_w\" -q dataout_w_cnt");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"dataout_w_ori_reg_en\" -d \"dataout_w_cnt_w\" -q dataout_w_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dataout_w_cnt <= {13{1'b0}};
   end else begin
       if ((dataout_w_cnt_reg_en) == 1'b1) begin
           dataout_w_cnt <= dataout_w_cnt_w;
       // VCS coverage off
       end else if ((dataout_w_cnt_reg_en) == 1'b0) begin
       end else begin
           dataout_w_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dataout_w_ori <= {13{1'b0}};
   end else begin
       if ((dataout_w_ori_reg_en) == 1'b1) begin
           dataout_w_ori <= dataout_w_cnt_w;
       // VCS coverage off
       end else if ((dataout_w_ori_reg_en) == 1'b0) begin
       end else begin
           dataout_w_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// input channel coordinate counter, only feature  //////////////////////////
assign {mon_datain_c_cnt_inc,datain_c_cnt_inc} = datain_c_cnt + 1'b1;
assign is_last_channel = (datain_c_cnt == datain_channel_cmp);
assign datain_c_cnt_w = layer_st ? 11'b0 : dl_channel_end ? 11'b0 : datain_c_cnt_inc;
assign datain_c_cnt_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_block_end);
//: &eperl::flop("-nodeclare   -rval \"{11{1'b0}}\"  -en \"datain_c_cnt_reg_en\" -d \"datain_c_cnt_w\" -q datain_c_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_c_cnt <= {11{1'b0}};
   end else begin
       if ((datain_c_cnt_reg_en) == 1'b1) begin
           datain_c_cnt <= datain_c_cnt_w;
       // VCS coverage off
       end else if ((datain_c_cnt_reg_en) == 1'b0) begin
       end else begin
           datain_c_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// input width coordinate counter, feature/image dedicated counter //////////////////////////
assign datain_w_cnt_st = (is_img) ? 14'b0 : (is_winograd) ? 14'h2 : 13'b0 - reg2dp_pad_left;
assign {mon_datain_w_cnt_inc,datain_w_cnt_inc} = (is_winograd_d1[3]) ? (datain_w_cnt + 2'h2) : (datain_w_cnt + conv_x_stride);
//full data cube w counter,start form negtive, only for feature data. non-image, by element
assign datain_w_cnt_w = layer_st ? datain_w_cnt_st :
                        (is_stripe_end & ~dl_channel_end) ? datain_w_ori :
                        is_w_end ? datain_w_cnt_st :
                        datain_w_cnt_inc;
assign dl_w_offset_ext = dl_w_offset * x_dilate;
assign {mon_datain_w_cur,datain_w_cur} = datain_w_cnt + dl_w_offset_ext; //by element
assign datain_w_cnt_reg_en = layer_st | (dat_exec_valid & is_batch_end & is_sub_h_end & ~is_img_d1[0]);
assign datain_w_ori_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_channel_end & ~is_img_d1[1]);
//notice:after sub_h T, pixel_x_add elements in W direction is used by CMAC
assign pixel_x_cnt_add = (is_sub_h_end) ? pixel_x_add : 6'b0;
//assign {mon_pixel_w_cnt_w,pixel_w_cnt_w} = (layer_st_d1) ? {{11{1'b0}}, pixel_x_init} :
// (is_stripe_end & dl_block_end & dl_channel_end & is_w_end) ? {{11{1'b0}}, pixel_x_init} :
// (is_stripe_end & dl_block_end & dl_channel_end & ~is_w_end) ? (pixel_w_ch_ori + pixel_ch_stride) :
// (is_stripe_end & dl_block_end & ~dl_channel_end) ? (pixel_w_ch_ori + pixel_x_init_offset) :
// (is_stripe_end & ~dl_block_end) ? {1'b0, pixel_w_ori} :
// (pixel_w_cnt + pixel_x_cnt_add);
//channel count.
wire [12:0] total_channel_op = (reg2dp_weight_channel_ext[6 -1:0]=={6{1'b0}}) ?
                        reg2dp_weight_channel_ext[12:6] : reg2dp_weight_channel_ext[12:6]+1'b1;
reg [12:0] channel_op_cnt;
wire mon_channel_op_cnt_nxt;
wire [12:0] channel_op_cnt_nxt;
assign {mon_channel_op_cnt_nxt, channel_op_cnt_nxt} = dl_channel_end&is_stripe_end ? 13'h2 :
                                                        dl_block_end&is_stripe_end ? channel_op_cnt + 1'b1 :
                                                        channel_op_cnt;
//: &eperl::flop("-q channel_op_cnt  -d \"channel_op_cnt_nxt\"  -wid 13  -rval \"13'h2\" -nodeclare ");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       channel_op_cnt <= 13'h2;
   end else begin
       channel_op_cnt <= channel_op_cnt_nxt;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
wire next_is_last_channel = (channel_op_cnt >= total_channel_op);
//notice, after pre-extention, image weight w_total <=128
assign {mon_pixel_w_cnt_w,pixel_w_cnt_w} = (layer_st_d1) ? {{11{1'b0}}, pixel_x_init} :
                        (is_stripe_end & dl_block_end & dl_channel_end & is_w_end) ? {{11{1'b0}}, pixel_x_init} :
                        (is_stripe_end & dl_block_end & dl_channel_end & ~is_w_end) ? (pixel_w_ch_ori + pixel_ch_stride) :
//(is_stripe_end & dl_block_end & ~dl_channel_end) ? (pixel_w_ori + dl_in_pd_d0[16:10]) :
                        (is_stripe_end & dl_block_end & next_is_last_channel) ? (pixel_w_ori + pixel_x_init_offset) :
                        (is_stripe_end & dl_block_end & ~next_is_last_channel) ? (pixel_w_ori + 8'h40  ) :
                        (is_stripe_end & ~dl_block_end) ? {1'b0, pixel_w_ori} :
                        (pixel_w_cnt + pixel_x_cnt_add);
assign pixel_w_cur = {{6 -1{1'b0}},pixel_w_cnt[15:6]}; //by entry 
assign pixel_w_cnt_reg_en = layer_st_d1 | (dat_exec_valid & is_img_d1[2] & (is_sub_h_end | is_w_end));
assign pixel_w_ori_reg_en = layer_st_d1 | (dat_exec_valid & is_img_d1[3] & is_stripe_end & dl_block_end);
assign pixel_ch_ori_reg_en = layer_st_d1 | (dat_exec_valid & is_img_d1[4] & is_stripe_end & dl_block_end & dl_channel_end);
assign pixel_force_fetch = (is_img_d1[0] & dat_req_stripe_st) ? 1'b1 : (pixel_force_clr_d1) ? 1'b0 : pixel_force_fetch_d1;
assign pixel_force_clr = is_img_d1[0] & is_sub_h_end & (pixel_force_fetch | pixel_force_fetch_d1);
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_w_cnt_reg_en\" -d \"datain_w_cnt_w\" -q datain_w_cnt");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_w_ori_reg_en\" -d \"datain_w_cnt_w\" -q datain_w_ori");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"pixel_w_cnt_reg_en\" -d \"pixel_w_cnt_w\" -q pixel_w_cnt");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"pixel_w_ori_reg_en\" -d \"pixel_w_cnt_w\" -q pixel_w_ori");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"pixel_ch_ori_reg_en\" -d \"pixel_w_cnt_w\" -q pixel_w_ch_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_w_cnt <= {14{1'b0}};
   end else begin
       if ((datain_w_cnt_reg_en) == 1'b1) begin
           datain_w_cnt <= datain_w_cnt_w;
       // VCS coverage off
       end else if ((datain_w_cnt_reg_en) == 1'b0) begin
       end else begin
           datain_w_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_w_ori <= {14{1'b0}};
   end else begin
       if ((datain_w_ori_reg_en) == 1'b1) begin
           datain_w_ori <= datain_w_cnt_w;
       // VCS coverage off
       end else if ((datain_w_ori_reg_en) == 1'b0) begin
       end else begin
           datain_w_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_w_cnt <= {16{1'b0}};
   end else begin
       if ((pixel_w_cnt_reg_en) == 1'b1) begin
           pixel_w_cnt <= pixel_w_cnt_w;
       // VCS coverage off
       end else if ((pixel_w_cnt_reg_en) == 1'b0) begin
       end else begin
           pixel_w_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_w_ori <= {16{1'b0}};
   end else begin
       if ((pixel_w_ori_reg_en) == 1'b1) begin
           pixel_w_ori <= pixel_w_cnt_w;
       // VCS coverage off
       end else if ((pixel_w_ori_reg_en) == 1'b0) begin
       end else begin
           pixel_w_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_w_ch_ori <= {16{1'b0}};
   end else begin
       if ((pixel_ch_ori_reg_en) == 1'b1) begin
           pixel_w_ch_ori <= pixel_w_cnt_w;
       // VCS coverage off
       end else if ((pixel_ch_ori_reg_en) == 1'b0) begin
       end else begin
           pixel_w_ch_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// input height coordinate counter, feature/image both  //////////////////////////
// full data cube h counter, start form negative
assign datain_h_cnt_st = (is_winograd) ? 14'b0 : 14'b0 - reg2dp_pad_top;
assign {mon_datain_h_cnt_inc, datain_h_cnt_inc} = datain_h_cnt + conv_y_stride;
assign datain_h_cnt_w = (layer_st | (is_stripe_end & dl_group_end)) ? datain_h_cnt_st :
                        (is_stripe_end & ~dl_channel_end) ? datain_h_ori :
                        is_w_end ? datain_h_cnt_inc :
                        datain_h_cnt;
assign datain_h_cnt_reg_en = layer_st | (dat_exec_valid & ((is_stripe_end & ~dl_channel_end) | is_w_end));
assign datain_h_ori_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_channel_end);
assign dl_h_offset_ext = dl_h_offset * y_dilate;
assign {mon_datain_h_cur,datain_h_cur} = datain_h_cnt + dl_h_offset_ext + sub_h_cnt;
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_h_cnt_reg_en\" -d \"datain_h_cnt_w\" -q datain_h_cnt");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_h_ori_reg_en\" -d \"datain_h_cnt_w\" -q datain_h_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_h_cnt <= {14{1'b0}};
   end else begin
       if ((datain_h_cnt_reg_en) == 1'b1) begin
           datain_h_cnt <= datain_h_cnt_w;
       // VCS coverage off
       end else if ((datain_h_cnt_reg_en) == 1'b0) begin
       end else begin
           datain_h_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_h_ori <= {14{1'b0}};
   end else begin
       if ((datain_h_ori_reg_en) == 1'b1) begin
           datain_h_ori <= datain_h_cnt_w;
       // VCS coverage off
       end else if ((datain_h_ori_reg_en) == 1'b0) begin
       end else begin
           datain_h_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// fetch valid generate //////////////////////////
assign dat_conv_req_dummy = (datain_w_cur[13 ]) | (datain_w_cur > {1'b0, datain_width_cmp})
                            | (datain_h_cur[13 ]) | (datain_h_cur > {1'b0, datain_height_cmp});
assign dat_wg_req_dummy = 1'b0;
assign dat_wg_req_skip = ((|datain_w_cur[13:2]) & datain_w_cur[1] & (|stripe_cnt[6:1]));
assign dat_img_req_dummy = (datain_h_cur[13]) | (datain_h_cur > {1'b0, datain_height_cmp});
//w address(in entry) is bigger than avilable entrys
assign dat_img_req_skip = ({{15 -12{1'b0}},w_bias_w[13:2]} > entries_cmp[15 -1:0]);
assign dat_req_dummy = is_img_d1[5] ? dat_img_req_dummy : is_winograd_d1[4] ? dat_wg_req_dummy : dat_conv_req_dummy;
assign dat_req_skip = (is_winograd_d1[5] & dat_wg_req_skip) | (is_img_d1[6] & dat_img_req_skip);
assign dat_req_valid = (dat_exec_valid & ~dat_req_dummy & ~dat_req_skip);
//Add corner case
assign dat_req_sub_c_w = ~is_img_d1[7] ? datain_c_cnt[0] : dl_block_end;
assign dat_req_sub_w_w = is_winograd_d1[6] ? {1'b0, ~datain_w_cur[1]} : datain_w_cur[1:0];
assign dat_req_sub_w_st_en = dat_exec_valid & (sub_h_cnt == 2'h0);
assign dat_req_batch_index = batch_cnt;
assign dat_req_stripe_st = dl_pvld;
assign dat_req_stripe_end = is_stripe_equal & dat_pipe_valid;
assign dat_req_channel_end = dl_channel_end;
assign dat_req_layer_end = dl_layer_end;
// PKT_PACK_WIRE( nvdla_stripe_info , dat_req_ , dat_req_flag_w )
assign dat_req_flag_w[4:0] = dat_req_batch_index[4:0];
assign dat_req_flag_w[5] = dat_req_stripe_st ;
assign dat_req_flag_w[6] = dat_req_stripe_end ;
assign dat_req_flag_w[7] = dat_req_channel_end ;
assign dat_req_flag_w[8] = dat_req_layer_end ;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_req_valid\" -q dat_req_valid_d1");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid\" -d \"dat_req_sub_w_w\" -q dat_req_sub_w_d1");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid\" -d \"sub_h_cnt\" -q dat_req_sub_h_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"dat_req_sub_c_w\" -q dat_req_sub_c_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"is_last_channel\" -q dat_req_ch_end_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"dat_req_dummy\" -q dat_req_dummy_d1");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid\" -d \"dl_cur_sub_h\" -q dat_req_cur_sub_h_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_req_sub_w_st_en\" -d \"dat_req_stripe_st\" -q dat_req_sub_w_st_d1");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_exec_valid\" -d \"dat_req_flag_w\" -q dat_req_flag_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"dl_dat_release & is_stripe_equal & dat_pipe_valid\" -q dat_req_rls_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"pixel_force_fetch\" -q pixel_force_fetch_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"pixel_force_clr\" -q pixel_force_clr_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_valid_d1 <= 1'b0;
   end else begin
       dat_req_valid_d1 <= dat_req_valid;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_d1 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_sub_w_d1 <= dat_req_sub_w_w;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_sub_w_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_d1 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_sub_h_d1 <= sub_h_cnt;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_sub_h_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_c_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_sub_c_d1 <= dat_req_sub_c_w;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_sub_c_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_ch_end_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_ch_end_d1 <= is_last_channel;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_ch_end_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_dummy_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_dummy_d1 <= dat_req_dummy;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_dummy_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_cur_sub_h_d1 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_cur_sub_h_d1 <= dl_cur_sub_h;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_cur_sub_h_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_st_d1 <= 1'b0;
   end else begin
       if ((dat_req_sub_w_st_en) == 1'b1) begin
           dat_req_sub_w_st_d1 <= dat_req_stripe_st;
       // VCS coverage off
       end else if ((dat_req_sub_w_st_en) == 1'b0) begin
       end else begin
           dat_req_sub_w_st_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_flag_d1 <= {9{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_flag_d1 <= dat_req_flag_w;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_flag_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_rls_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_rls_d1 <= dl_dat_release & is_stripe_equal & dat_pipe_valid;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_rls_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_force_fetch_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           pixel_force_fetch_d1 <= pixel_force_fetch;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           pixel_force_fetch_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_force_clr_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           pixel_force_clr_d1 <= pixel_force_clr;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           pixel_force_clr_d1 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// generate data read address                         /////
//////////////////////////////////////////////////////////////
////////////////////////// data read index generator: 1st stage //////////////////////////
//channel bias, by w_in element
//assign c_bias_add = (~is_img_d1[8] & datain_c_cnt[0]) ? datain_width[12 -1:0] : 12'b0;
assign c_bias_add = (~is_img_d1[8]) ? datain_width[12 -1:0] : 12'b0;
assign {mon_c_bias_w, c_bias_w} = layer_st ? 13'b0 : (is_stripe_end & dl_channel_end) ? 13'b0 : c_bias + c_bias_add;
assign c_bias_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_block_end);
assign c_bias_d1_reg_en = (c_bias != c_bias_d1);
//height bias, by element
assign {mon_h_bias_0_w,h_bias_0_w} = datain_h_cnt[13:0] * h_bias_0_stride;
assign {mon_h_bias_1_w,h_bias_1_w} = dl_h_offset * h_bias_1_stride;
assign {mon_h_bias_2_w,h_bias_2_w} = batch_cnt * h_bias_2_stride;
assign {mon_h_bias_3_w,h_bias_3_w} = layer_st ? 13'b0 :sub_h_cnt * h_bias_3_stride;
assign h_bias_reg_en[0] = dat_exec_valid;
assign h_bias_reg_en[1] = layer_st | (dat_exec_valid & (is_winograd_d1[7] | is_img_d1[9]));
//width bias, by entry in image, by element in feature data

assign w_bias_int8 = is_img_d1[10] ? {pixel_w_cur} : //by entry in image 
                     is_winograd_d1[8] ? {1'b0, datain_w_cnt} :
                     (~is_last_channel | is_winograd_d1[8]) ? {2'b0,datain_w_cur[12:0]} ://not last channel, by element
                     (dat_req_bytes > 8'h20) ? {2'b0,datain_w_cur[12:0]} : //last channel & request >1/2*entry
                     {3'b0, datain_w_cur[12:1]}; //last channel & request<=1/2*entry

assign w_bias_int8 = is_img_d1[10] ? {pixel_w_cur} : //by entry in image 
                     is_winograd_d1[8] ? {1'b0, datain_w_cnt} :
                     (~is_last_channel | is_winograd_d1[8]) ? {2'b0,datain_w_cur[12:0]} ://not last channel, by element
                     (dat_req_bytes > 8'h20) ? {2'b0,datain_w_cur[12:0]} : //last channel & request >1/2*entry
                     (dat_req_bytes <= 8'h10) ? {4'b0, datain_w_cur[12:2]} : //last channel & request <=1/4*entry
                     {3'b0, datain_w_cur[12:1]}; //last channel & (1/4*entry<request<=1/2*entry)
assign w_bias_w = w_bias_int8[13:0];
assign w_bias_reg_en = dat_exec_valid;
assign dat_req_base_d1 = dat_entry_st[13 -1:0];
//: my $kk=13;
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"c_bias_reg_en\" -d \"c_bias_w\" -q c_bias");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"c_bias_d1_reg_en\" -d \"c_bias\" -q c_bias_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[0]\" -d \"h_bias_0_w\" -q h_bias_0_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[0]\" -d \"h_bias_1_w\" -q h_bias_1_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[0]\" -d \"h_bias_2_w\" -q h_bias_2_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[1]\" -d \"h_bias_3_w\" -q h_bias_3_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"w_bias_reg_en\" -d \"w_bias_w\" -q w_bias_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       c_bias <= {13{1'b0}};
   end else begin
       if ((c_bias_reg_en) == 1'b1) begin
           c_bias <= c_bias_w;
       // VCS coverage off
       end else if ((c_bias_reg_en) == 1'b0) begin
       end else begin
           c_bias <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       c_bias_d1 <= {13{1'b0}};
   end else begin
       if ((c_bias_d1_reg_en) == 1'b1) begin
           c_bias_d1 <= c_bias;
       // VCS coverage off
       end else if ((c_bias_d1_reg_en) == 1'b0) begin
       end else begin
           c_bias_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_0_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[0]) == 1'b1) begin
           h_bias_0_d1 <= h_bias_0_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[0]) == 1'b0) begin
       end else begin
           h_bias_0_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_1_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[0]) == 1'b1) begin
           h_bias_1_d1 <= h_bias_1_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[0]) == 1'b0) begin
       end else begin
           h_bias_1_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_2_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[0]) == 1'b1) begin
           h_bias_2_d1 <= h_bias_2_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[0]) == 1'b0) begin
       end else begin
           h_bias_2_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_3_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[1]) == 1'b1) begin
           h_bias_3_d1 <= h_bias_3_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[1]) == 1'b0) begin
       end else begin
           h_bias_3_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       w_bias_d1 <= {13{1'b0}};
   end else begin
       if ((w_bias_reg_en) == 1'b1) begin
           w_bias_d1 <= w_bias_w;
       // VCS coverage off
       end else if ((w_bias_reg_en) == 1'b0) begin
       end else begin
           w_bias_d1 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// data read index generator: 2st stage //////////////////////////
wire [13 -1:0] dat_req_addr_minus1;
wire mon_dat_req_addr_minus1;
wire is_dat_req_addr_minus1_wrap;
wire [13 -1:0] dat_req_addr_minus1_wrap;
wire [13 -1:0] dat_req_addr_minus1_real;
assign {mon_h_bias_d1,h_bias_d1} = h_bias_0_d1 + h_bias_1_d1 + h_bias_2_d1 + h_bias_3_d1;
//assign {mon_dat_req_addr_sum,dat_req_addr_sum} = dat_req_base_d1 + c_bias_d1 + h_bias_d1 + w_bias_d1; //by entry
assign dat_req_addr_sum = dat_req_base_d1 + c_bias_d1 + h_bias_d1 + w_bias_d1; //by entry
assign is_dat_req_addr_wrap = (dat_req_addr_sum >= {1'b0,data_bank, {9{1'b0}}});
assign {mon_dat_req_addr_wrap,dat_req_addr_wrap} = dat_req_addr_sum[13:0] - {1'b0,data_bank, {9{1'b0}}};
assign dat_req_addr_w = (layer_st | dat_req_dummy_d1) ? {13{1'b1}} : is_dat_req_addr_wrap ? dat_req_addr_wrap : dat_req_addr_sum[13 -1:0]; //get the adress sends to cbuf
assign {mon_dat_req_addr_minus1,dat_req_addr_minus1} = dat_req_addr_w-1'b1;
assign is_dat_req_addr_minus1_wrap = (dat_req_addr_minus1 >= {data_bank, {9{1'b0}}}); //only one case: 0-1=ffff would introduce wrap  
assign dat_req_addr_minus1_wrap = {data_bank, {9{1'b1}}};
assign dat_req_addr_minus1_real = is_dat_req_addr_minus1_wrap ? dat_req_addr_minus1_wrap : dat_req_addr_minus1;
assign sc2buf_dat_rd_en_w = dat_req_valid_d1 & ((dat_req_addr_last != dat_req_addr_w) | pixel_force_fetch_d1);
assign dat_req_addr_last = (dat_req_sub_h_d1 == 2'h0) ? dat_req_sub_h_0_addr :
                           (dat_req_sub_h_d1 == 2'h1) ? dat_req_sub_h_1_addr :
                           (dat_req_sub_h_d1 == 2'h2) ? dat_req_sub_h_2_addr :
                           dat_req_sub_h_3_addr;
assign dat_req_sub_h_0_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h0));
assign dat_req_sub_h_1_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h1));
assign dat_req_sub_h_2_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h2));
assign dat_req_sub_h_3_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h3));

wire [13 -1:0] sc2buf_dat_rd_addr_w;
assign sc2buf_dat_rd_addr_w = dat_req_addr_w;
//: my $kk=13;
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_0_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_0_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_1_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_1_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_2_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_2_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_3_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_3_addr");
//: my $kk=13;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"sc2buf_dat_rd_en_w\" -q sc2buf_dat_rd_en");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"layer_st | sc2buf_dat_rd_en_w\" -d \"sc2buf_dat_rd_addr_w\" -q sc2buf_dat_rd_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"layer_st | sc2buf_dat_rd_en_w\" -d \"sc2buf_dat_rd_next1_addr_w\" -q sc2buf_dat_rd_next1_addr");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_pipe_valid_d1\" -q dat_pipe_valid_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_exec_valid_d1\" -q dat_exec_valid_d2");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_w_d1\" -q dat_req_sub_w_d2");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_h_d1\" -q dat_req_sub_h_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_c_d1\" -q dat_req_sub_c_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_ch_end_d1\" -q dat_req_ch_end_d2");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_bytes_d1\" -q dat_req_bytes_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_dummy_d1\" -q dat_req_dummy_d2");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_cur_sub_h_d1\" -q dat_req_cur_sub_h_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_w_st_d1\" -q dat_req_sub_w_st_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_rls_d1\" -q dat_req_rls_d2");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_flag_d1\" -q dat_req_flag_d2");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_0_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_0_addr_en) == 1'b1) begin
           dat_req_sub_h_0_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_0_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_0_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_1_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_1_addr_en) == 1'b1) begin
           dat_req_sub_h_1_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_1_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_1_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_2_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_2_addr_en) == 1'b1) begin
           dat_req_sub_h_2_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_2_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_2_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_3_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_3_addr_en) == 1'b1) begin
           dat_req_sub_h_3_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_3_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_3_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2buf_dat_rd_en <= 1'b0;
   end else begin
       sc2buf_dat_rd_en <= sc2buf_dat_rd_en_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2buf_dat_rd_addr <= {13{1'b1}};
   end else begin
       if ((layer_st | sc2buf_dat_rd_en_w) == 1'b1) begin
           sc2buf_dat_rd_addr <= sc2buf_dat_rd_addr_w;
       // VCS coverage off
       end else if ((layer_st | sc2buf_dat_rd_en_w) == 1'b0) begin
       end else begin
           sc2buf_dat_rd_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_pipe_valid_d2 <= 1'b0;
   end else begin
       dat_pipe_valid_d2 <= dat_pipe_valid_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_exec_valid_d2 <= 1'b0;
   end else begin
       dat_exec_valid_d2 <= dat_exec_valid_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_d2 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_w_d2 <= dat_req_sub_w_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_w_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_d2 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_h_d2 <= dat_req_sub_h_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_h_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_c_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_c_d2 <= dat_req_sub_c_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_c_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_ch_end_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_ch_end_d2 <= dat_req_ch_end_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_ch_end_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_bytes_d2 <= {8{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_bytes_d2 <= dat_req_bytes_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_bytes_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_dummy_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_dummy_d2 <= dat_req_dummy_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_dummy_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_cur_sub_h_d2 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_cur_sub_h_d2 <= dat_req_cur_sub_h_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_cur_sub_h_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_st_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_w_st_d2 <= dat_req_sub_w_st_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_w_st_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_rls_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_rls_d2 <= dat_req_rls_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_rls_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_flag_d2 <= {9{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_flag_d2 <= dat_req_flag_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_flag_d2 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// sideband pipeline                                  /////
//////////////////////////////////////////////////////////////
assign dat_req_pipe_pvld = dat_pipe_valid_d2;
assign dat_req_pipe_sub_w = dat_req_sub_w_d2;
assign dat_req_pipe_sub_h = dat_req_sub_h_d2;
assign dat_req_pipe_sub_c = dat_req_sub_c_d2;
assign dat_req_pipe_ch_end = dat_req_ch_end_d2;
assign dat_req_pipe_bytes = dat_req_bytes_d2;
assign dat_req_pipe_dummy = dat_req_dummy_d2;
assign dat_req_pipe_cur_sub_h = dat_req_cur_sub_h_d2;
assign dat_req_pipe_sub_w_st = dat_req_sub_w_st_d2;
assign dat_req_pipe_rls = dat_req_rls_d2;
assign dat_req_pipe_flag = dat_req_flag_d2;
assign dat_req_exec_pvld = dat_exec_valid_d2;
assign dat_req_exec_dummy = dat_req_dummy_d2;
assign dat_req_exec_sub_h = dat_req_sub_h_d2;
// PKT_PACK_WIRE( csc_dat_req_pkg , dat_req_pipe_ , dat_req_pipe_pd )
assign dat_req_pipe_pd[1:0] = dat_req_pipe_sub_w[1:0];
assign dat_req_pipe_pd[3:2] = dat_req_pipe_sub_h[1:0];
assign dat_req_pipe_pd[4] = dat_req_pipe_sub_c ;
assign dat_req_pipe_pd[5] = dat_req_pipe_ch_end ;
assign dat_req_pipe_pd[6] = 1'b0 ;
assign dat_req_pipe_pd[14:7] = dat_req_pipe_bytes[7:0];
assign dat_req_pipe_pd[16:15] = dat_req_pipe_cur_sub_h[1:0];
assign dat_req_pipe_pd[17] = dat_req_pipe_dummy ;
assign dat_req_pipe_pd[18] = dat_req_pipe_sub_w_st ;
assign dat_req_pipe_pd[19] = dat_req_pipe_rls ;
assign dat_req_pipe_pd[28:20] = dat_req_pipe_flag[8:0];
//add latency for data request contorl signal
//: my $pipe_depth = 6;
//: my $i;
//: my $j;
//: if($pipe_depth == 0) {
//: print "assign dat_rsp_pipe_pvld = dat_req_pipe_pvld;\n";
//: print "assign dat_rsp_pipe_pd = dat_req_pipe_pd;\n";
//: print "assign dat_rsp_exec_pvld = dat_req_exec_pvld;\n";
//: print "assign dat_rsp_exec_dummy = dat_req_exec_dummy;\n";
//: print "assign dat_rsp_exec_sub_h = dat_req_exec_sub_h;\n\n";
//: } else {
//: print "assign dat_rsp_pipe_pvld_d0 = dat_req_pipe_pvld;\n";
//: print "assign dat_rsp_pipe_pd_d0 = dat_req_pipe_pd;\n";
//: print "assign dat_rsp_exec_pvld_d0 = dat_req_exec_pvld;\n";
//: print "assign dat_rsp_exec_dummy_d0 = dat_req_exec_dummy;\n";
//: print "assign dat_rsp_exec_sub_h_d0 = dat_req_exec_sub_h;\n\n";
//: for($i = 0; $i < $pipe_depth; $i ++) {
//: $j = $i + 1;
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -d \"dat_rsp_pipe_pvld_d${i}\"  -q dat_rsp_pipe_pvld_d${j}");
//: &eperl::flop("-wid 29  -rval \"{29{1'b0}}\" -en \"dat_rsp_pipe_pvld_d${i}\" -d \"dat_rsp_pipe_pd_d${i}\"    -q dat_rsp_pipe_pd_d${j}");
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -d \"dat_rsp_exec_pvld_d${i}\"  -q dat_rsp_exec_pvld_d${j}");
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -en \"dat_rsp_exec_pvld_d${i}\" -d \"dat_rsp_exec_dummy_d${i}\" -q dat_rsp_exec_dummy_d${j}");
//: &eperl::flop("-wid 2   -rval \"{2{1'b0}}\"  -en \"dat_rsp_exec_pvld_d${i}\" -d \"dat_rsp_exec_sub_h_d${i}\" -q dat_rsp_exec_sub_h_d${j}");
//: }
//: print "assign dat_rsp_pipe_pvld = dat_rsp_pipe_pvld_d${i};\n";
//: print "assign dat_rsp_pipe_pd = dat_rsp_pipe_pd_d${i};\n";
//: print "assign dat_rsp_exec_pvld = dat_rsp_exec_pvld_d${i};\n";
//: print "assign dat_rsp_exec_dummy = dat_rsp_exec_dummy_d${i};\n";
//: print "assign dat_rsp_exec_sub_h = dat_rsp_exec_sub_h_d${i};\n\n";
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_rsp_pipe_pvld_d0 = dat_req_pipe_pvld;
assign dat_rsp_pipe_pd_d0 = dat_req_pipe_pd;
assign dat_rsp_exec_pvld_d0 = dat_req_exec_pvld;
assign dat_rsp_exec_dummy_d0 = dat_req_exec_dummy;
assign dat_rsp_exec_sub_h_d0 = dat_req_exec_sub_h;

reg  dat_rsp_pipe_pvld_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d1 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d1 <= dat_rsp_pipe_pvld_d0;
   end
end
reg [28:0] dat_rsp_pipe_pd_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d1 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d0) == 1'b1) begin
           dat_rsp_pipe_pd_d1 <= dat_rsp_pipe_pd_d0;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d1 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d1 <= dat_rsp_exec_pvld_d0;
   end
end
reg  dat_rsp_exec_dummy_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d1 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d0) == 1'b1) begin
           dat_rsp_exec_dummy_d1 <= dat_rsp_exec_dummy_d0;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d1 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d0) == 1'b1) begin
           dat_rsp_exec_sub_h_d1 <= dat_rsp_exec_sub_h_d0;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d2 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d2 <= dat_rsp_pipe_pvld_d1;
   end
end
reg [28:0] dat_rsp_pipe_pd_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d2 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d1) == 1'b1) begin
           dat_rsp_pipe_pd_d2 <= dat_rsp_pipe_pd_d1;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d2 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d2 <= dat_rsp_exec_pvld_d1;
   end
end
reg  dat_rsp_exec_dummy_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d2 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d1) == 1'b1) begin
           dat_rsp_exec_dummy_d2 <= dat_rsp_exec_dummy_d1;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d2 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d1) == 1'b1) begin
           dat_rsp_exec_sub_h_d2 <= dat_rsp_exec_sub_h_d1;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d3 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d3 <= dat_rsp_pipe_pvld_d2;
   end
end
reg [28:0] dat_rsp_pipe_pd_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d3 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d2) == 1'b1) begin
           dat_rsp_pipe_pd_d3 <= dat_rsp_pipe_pd_d2;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d3 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d3 <= dat_rsp_exec_pvld_d2;
   end
end
reg  dat_rsp_exec_dummy_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d3 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d2) == 1'b1) begin
           dat_rsp_exec_dummy_d3 <= dat_rsp_exec_dummy_d2;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d3 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d2) == 1'b1) begin
           dat_rsp_exec_sub_h_d3 <= dat_rsp_exec_sub_h_d2;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d4 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d4 <= dat_rsp_pipe_pvld_d3;
   end
end
reg [28:0] dat_rsp_pipe_pd_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d4 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d3) == 1'b1) begin
           dat_rsp_pipe_pd_d4 <= dat_rsp_pipe_pd_d3;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d4 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d4 <= dat_rsp_exec_pvld_d3;
   end
end
reg  dat_rsp_exec_dummy_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d4 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d3) == 1'b1) begin
           dat_rsp_exec_dummy_d4 <= dat_rsp_exec_dummy_d3;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d4 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d3) == 1'b1) begin
           dat_rsp_exec_sub_h_d4 <= dat_rsp_exec_sub_h_d3;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d5 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d5 <= dat_rsp_pipe_pvld_d4;
   end
end
reg [28:0] dat_rsp_pipe_pd_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d5 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d4) == 1'b1) begin
           dat_rsp_pipe_pd_d5 <= dat_rsp_pipe_pd_d4;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d4) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d5 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d5 <= dat_rsp_exec_pvld_d4;
   end
end
reg  dat_rsp_exec_dummy_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d5 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d4) == 1'b1) begin
           dat_rsp_exec_dummy_d5 <= dat_rsp_exec_dummy_d4;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d4) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d5 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d4) == 1'b1) begin
           dat_rsp_exec_sub_h_d5 <= dat_rsp_exec_sub_h_d4;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d4) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d6 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d6 <= dat_rsp_pipe_pvld_d5;
   end
end
reg [28:0] dat_rsp_pipe_pd_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d6 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d5) == 1'b1) begin
           dat_rsp_pipe_pd_d6 <= dat_rsp_pipe_pd_d5;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d5) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d6 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d6 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d6 <= dat_rsp_exec_pvld_d5;
   end
end
reg  dat_rsp_exec_dummy_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d6 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d5) == 1'b1) begin
           dat_rsp_exec_dummy_d6 <= dat_rsp_exec_dummy_d5;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d5) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d6 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d6 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d5) == 1'b1) begin
           dat_rsp_exec_sub_h_d6 <= dat_rsp_exec_sub_h_d5;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d5) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d6 <= 'bx;
       // VCS coverage on
       end
   end
end
assign dat_rsp_pipe_pvld = dat_rsp_pipe_pvld_d6;
assign dat_rsp_pipe_pd = dat_rsp_pipe_pd_d6;
assign dat_rsp_exec_pvld = dat_rsp_exec_pvld_d6;
assign dat_rsp_exec_dummy = dat_rsp_exec_dummy_d6;
assign dat_rsp_exec_sub_h = dat_rsp_exec_sub_h_d6;


//| eperl: generated_end (DO NOT EDIT ABOVE)
// PKT_UNPACK_WIRE( csc_dat_req_pkg , dat_rsp_pipe_ , dat_rsp_pipe_pd )
assign dat_rsp_pipe_sub_w[1:0] = dat_rsp_pipe_pd[1:0];
assign dat_rsp_pipe_sub_h[1:0] = dat_rsp_pipe_pd[3:2];
assign dat_rsp_pipe_sub_c = dat_rsp_pipe_pd[4];
assign dat_rsp_pipe_ch_end = dat_rsp_pipe_pd[5];
assign dat_rsp_pipe_bytes[7:0] = dat_rsp_pipe_pd[14:7];
assign dat_rsp_pipe_cur_sub_h[1:0] = dat_rsp_pipe_pd[16:15];
assign dat_rsp_pipe_dummy = dat_rsp_pipe_pd[17];
assign dat_rsp_pipe_sub_w_st = dat_rsp_pipe_pd[18];
assign dat_rsp_pipe_rls = dat_rsp_pipe_pd[19];
assign dat_rsp_pipe_flag[8:0] = dat_rsp_pipe_pd[28:20];
//////////////////////////////////////////////////////////////
///// dl data cache                                      /////
//////////////////////////////////////////////////////////////
assign dat_l0c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h0));
assign dat_l1c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h1));
assign dat_l2c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h2));
assign dat_l3c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h3));
//only winograd/image
assign dat_l0c1_en = (dat_wg_adv & ~dat_rsp_exec_sub_h[0]) | (is_img_d1[12] & dat_l0c0_en & ~dat_l0c0_dummy);
assign dat_l1c1_en = (dat_wg_adv & dat_rsp_exec_sub_h[0]) | (is_img_d1[13] & dat_l1c0_en & ~dat_l1c0_dummy);
assign dat_l2c1_en = (is_img_d1[15] & dat_l2c0_en & ~dat_l2c0_dummy);
assign dat_l3c1_en = (is_img_d1[16] & dat_l3c0_en & ~dat_l3c0_dummy);
assign dat_dummy_l0_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h0);
assign dat_dummy_l1_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h1);
assign dat_dummy_l2_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h2);
assign dat_dummy_l3_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h3);
assign dat_wg_adv = sc2buf_dat_rd_valid & is_winograd_d1[11] & ~dat_rsp_pipe_sub_w_st;
assign dat_l0c0_dummy_w = dat_l0c0_en ? 1'b0 : dat_dummy_l0_en ? 1'b1 : dat_l0c0_dummy;
assign dat_l1c0_dummy_w = dat_l1c0_en ? 1'b0 : dat_dummy_l1_en ? 1'b1 : dat_l1c0_dummy;
assign dat_l2c0_dummy_w = dat_l2c0_en ? 1'b0 : dat_dummy_l2_en ? 1'b1 : dat_l2c0_dummy;
assign dat_l3c0_dummy_w = dat_l3c0_en ? 1'b0 : dat_dummy_l3_en ? 1'b1 : dat_l3c0_dummy;
assign dat_l0c1_dummy_w = dat_l0c1_en ? 1'b0 : (dat_l0_set) ? dat_l0c0_dummy : dat_l0c1_dummy;
assign dat_l1c1_dummy_w = dat_l1c1_en ? 1'b0 : (dat_l1_set & (|sub_h_total_g2)) ? dat_l1c0_dummy : dat_l1c1_dummy;
assign dat_l2c1_dummy_w = dat_l2c1_en ? 1'b0 : (dat_l2_set & sub_h_total_g2[1]) ? dat_l2c0_dummy : dat_l2c1_dummy;
assign dat_l3c1_dummy_w = dat_l3c1_en ? 1'b0 : (dat_l3_set & sub_h_total_g2[1]) ? dat_l3c0_dummy : dat_l3c1_dummy;
assign dat_l0_set = dat_l0c0_en | dat_dummy_l0_en;
assign dat_l1_set = dat_l1c0_en | dat_dummy_l1_en;
assign dat_l2_set = dat_l2c0_en | dat_dummy_l2_en;
assign dat_l3_set = dat_l3c0_en | dat_dummy_l3_en;
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l0c0_dummy_w\" -q dat_l0c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l1c0_dummy_w\" -q dat_l1c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l2c0_dummy_w\" -q dat_l2c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l3c0_dummy_w\" -q dat_l3c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l0c1_dummy_w\" -q dat_l0c1_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l1c1_dummy_w\" -q dat_l1c1_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l2c1_dummy_w\" -q dat_l2c1_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l3c1_dummy_w\" -q dat_l3c1_dummy");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l0c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l0c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l1c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l1c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l2c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l2c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l3c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l3c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l0c1_en\" -d dat_l0c0 -q dat_l0c1 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l1c1_en\" -d dat_l1c0 -q dat_l1c1 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l2c1_en\" -d dat_l2c0 -q dat_l2c1 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l3c1_en\" -d dat_l3c0 -q dat_l3c1 ");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l0c0_dummy <= 1'b1;
   end else begin
       dat_l0c0_dummy <= dat_l0c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l1c0_dummy <= 1'b1;
   end else begin
       dat_l1c0_dummy <= dat_l1c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l2c0_dummy <= 1'b1;
   end else begin
       dat_l2c0_dummy <= dat_l2c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l3c0_dummy <= 1'b1;
   end else begin
       dat_l3c0_dummy <= dat_l3c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l0c1_dummy <= 1'b1;
   end else begin
       dat_l0c1_dummy <= dat_l0c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l1c1_dummy <= 1'b1;
   end else begin
       dat_l1c1_dummy <= dat_l1c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l2c1_dummy <= 1'b1;
   end else begin
       dat_l2c1_dummy <= dat_l2c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l3c1_dummy <= 1'b1;
   end else begin
       dat_l3c1_dummy <= dat_l3c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l0c0_en) == 1'b1) begin
           dat_l0c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l0c0_en) == 1'b0) begin
       end else begin
           dat_l0c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l1c0_en) == 1'b1) begin
           dat_l1c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l1c0_en) == 1'b0) begin
       end else begin
           dat_l1c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l2c0_en) == 1'b1) begin
           dat_l2c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l2c0_en) == 1'b0) begin
       end else begin
           dat_l2c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l3c0_en) == 1'b1) begin
           dat_l3c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l3c0_en) == 1'b0) begin
       end else begin
           dat_l3c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l0c1_en) == 1'b1) begin
           dat_l0c1 <= dat_l0c0;
       // VCS coverage off
       end else if ((dat_l0c1_en) == 1'b0) begin
       end else begin
           dat_l0c1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l1c1_en) == 1'b1) begin
           dat_l1c1 <= dat_l1c0;
       // VCS coverage off
       end else if ((dat_l1c1_en) == 1'b0) begin
       end else begin
           dat_l1c1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l2c1_en) == 1'b1) begin
           dat_l2c1 <= dat_l2c0;
       // VCS coverage off
       end else if ((dat_l2c1_en) == 1'b0) begin
       end else begin
           dat_l2c1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l3c1_en) == 1'b1) begin
           dat_l3c1 <= dat_l3c0;
       // VCS coverage off
       end else if ((dat_l3c1_en) == 1'b0) begin
       end else begin
           dat_l3c1 <= 'bx;
       // VCS coverage on
       end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// response contorl                                   /////
//////////////////////////////////////////////////////////////
// PKT_PACK_WIRE( csc_dat_rsp_pkg , dat_rsp_pipe_ , dat_rsp_pd_d0 )
assign dat_rsp_pd_d0[1:0] = dat_rsp_pipe_sub_w[1:0];
assign dat_rsp_pd_d0[3:2] = dat_rsp_pipe_sub_h[1:0];
assign dat_rsp_pd_d0[4] = dat_rsp_pipe_sub_c ;
assign dat_rsp_pd_d0[5] = dat_rsp_pipe_ch_end ;
assign dat_rsp_pd_d0[6] = 1'b0 ;
assign dat_rsp_pd_d0[14:7] = dat_rsp_pipe_bytes[7:0];
assign dat_rsp_pd_d0[16:15] = dat_rsp_pipe_cur_sub_h[1:0];
assign dat_rsp_pd_d0[17] = dat_rsp_pipe_rls ;
assign dat_rsp_pd_d0[26:18] = dat_rsp_pipe_flag[8:0];
//add latency
//: my $delay_depth = 4;
//: my $i;
//: my $j;
//:
//: print "assign dat_rsp_pvld_d0 = dat_rsp_pipe_pvld;\n";
//: for($i = 0; $i < $delay_depth; $i ++) {
//: $j = $i + 1;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"           -d \"dat_rsp_pvld_d${i}\"   -q dat_rsp_pvld_d${j}");
//: &eperl::flop("-nodeclare   -rval \"{27{1'b0}}\"     -en \"dat_rsp_pvld_d${i}\"  -d \"dat_rsp_pd_d${i}\" -q dat_rsp_pd_d${j}");
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_rsp_pvld_d0 = dat_rsp_pipe_pvld;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d1 <= 1'b0;
   end else begin
       dat_rsp_pvld_d1 <= dat_rsp_pvld_d0;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d1 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d0) == 1'b1) begin
           dat_rsp_pd_d1 <= dat_rsp_pd_d0;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d2 <= 1'b0;
   end else begin
       dat_rsp_pvld_d2 <= dat_rsp_pvld_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d2 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d1) == 1'b1) begin
           dat_rsp_pd_d2 <= dat_rsp_pd_d1;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d3 <= 1'b0;
   end else begin
       dat_rsp_pvld_d3 <= dat_rsp_pvld_d2;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d3 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d2) == 1'b1) begin
           dat_rsp_pd_d3 <= dat_rsp_pd_d2;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d4 <= 1'b0;
   end else begin
       dat_rsp_pvld_d4 <= dat_rsp_pvld_d3;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d4 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d3) == 1'b1) begin
           dat_rsp_pd_d4 <= dat_rsp_pd_d3;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dat_rsp_pvld = (sub_h_total_g3[2] & dat_rsp_pvld_d4) |
                      (sub_h_total_g3[1] & dat_rsp_pvld_d2) |
                      (sub_h_total_g3[0] & dat_rsp_pvld_d1);
assign dat_rsp_l0_pvld = dat_rsp_pvld_d1;
assign dat_rsp_l1_pvld = dat_rsp_pvld_d2;
assign dat_rsp_l2_pvld = dat_rsp_pvld_d3;
assign dat_rsp_l3_pvld = dat_rsp_pvld_d4;
assign dat_rsp_pd = ({27 {sub_h_total_g4[2]}} & dat_rsp_pd_d4) |
                    ({27 {sub_h_total_g4[1]}} & dat_rsp_pd_d2) |
                    ({27 {sub_h_total_g4[0]}} & dat_rsp_pd_d1);
assign dat_rsp_l0_sub_c = dat_rsp_pd_d1[4:4];
assign dat_rsp_l1_sub_c = dat_rsp_pd_d2[4:4];
assign dat_rsp_l2_sub_c = dat_rsp_pd_d3[4:4];
assign dat_rsp_l3_sub_c = dat_rsp_pd_d4[4:4];
assign dat_rsp_l0_flag = dat_rsp_pd_d1[26:18];
assign dat_rsp_l1_flag = dat_rsp_pd_d2[26:18];
assign dat_rsp_l2_flag = dat_rsp_pd_d3[26:18];
assign dat_rsp_l3_flag = dat_rsp_pd_d4[26:18];
assign dat_rsp_l0_stripe_end = dat_rsp_l0_flag[6:6];
assign dat_rsp_l1_stripe_end = dat_rsp_l1_flag[6:6];
assign dat_rsp_l2_stripe_end = dat_rsp_l2_flag[6:6];
assign dat_rsp_l3_stripe_end = dat_rsp_l3_flag[6:6];
// PKT_UNPACK_WIRE( csc_dat_rsp_pkg , dat_rsp_ , dat_rsp_pd )
assign dat_rsp_sub_w[1:0] = dat_rsp_pd[1:0];
assign dat_rsp_sub_h[1:0] = dat_rsp_pd[3:2];
assign dat_rsp_sub_c = dat_rsp_pd[4];
assign dat_rsp_ch_end = dat_rsp_pd[5];
assign dat_rsp_bytes[7:0] = dat_rsp_pd[14:7];
assign dat_rsp_cur_sub_h[1:0] = dat_rsp_pd[16:15];
assign dat_rsp_rls = dat_rsp_pd[17];
assign dat_rsp_flag[8:0] = dat_rsp_pd[26:18];
// PKT_UNPACK_WIRE( nvdla_stripe_info , dat_rsp_ , dat_rsp_flag )
assign dat_rsp_batch_index[4:0] = dat_rsp_flag[4:0];
assign dat_rsp_stripe_st = dat_rsp_flag[5];
assign dat_rsp_stripe_end = dat_rsp_flag[6];
assign dat_rsp_channel_end = dat_rsp_flag[7];
assign dat_rsp_layer_end = dat_rsp_flag[8];
assign rsp_sft_cnt_l0_sub = dat_l0c0_en ? 8'h40   : 8'h0;
assign rsp_sft_cnt_l1_sub = dat_l1c0_en ? 8'h40   : 8'h0;
assign rsp_sft_cnt_l2_sub = dat_l2c0_en ? 8'h40   : 8'h0;
assign rsp_sft_cnt_l3_sub = dat_l3c0_en ? 8'h40   : 8'h0;
////: &eperl::retime("-O stripe_begin_disable_jump_7T -i stripe_begin_disable_jump -stage 8 -clk nvdla_core_clk");
////: &eperl::flop("-q stripe_begin_disable_jump_8T -d stripe_begin_disable_jump_7T -clk nvdla_core_clk");
assign {mon_rsp_sft_cnt_l0_w,rsp_sft_cnt_l0_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l0 + pixel_x_byte_stride - rsp_sft_cnt_l0_sub);
assign {mon_rsp_sft_cnt_l1_w,rsp_sft_cnt_l1_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l1 + pixel_x_byte_stride - rsp_sft_cnt_l1_sub);
assign {mon_rsp_sft_cnt_l2_w,rsp_sft_cnt_l2_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l2 + pixel_x_byte_stride - rsp_sft_cnt_l2_sub);
assign {mon_rsp_sft_cnt_l3_w,rsp_sft_cnt_l3_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l3 + pixel_x_byte_stride - rsp_sft_cnt_l3_sub);
//the data frm cbuf's low Bytes is always needed. High Bytes maybe unneeded.
assign dat_rsp_l0_block_end = dat_rsp_l0_sub_c;
assign dat_rsp_l1_block_end = dat_rsp_l1_sub_c;
assign dat_rsp_l2_block_end = dat_rsp_l2_sub_c;
assign dat_rsp_l3_block_end = dat_rsp_l3_sub_c;
assign rsp_sft_cnt_l0_w = (layer_st) ? 8'h40   : //begin from C0
                          (dat_rsp_l0_stripe_end & ~dat_rsp_l0_block_end) ? rsp_sft_cnt_l0_ori :
                          (dat_rsp_l0_stripe_end & dat_rsp_l0_block_end) ? 8'h40   :
                          (dat_dummy_l0_en) ? (rsp_sft_cnt_l0_inc & 8'h3f) :
                          rsp_sft_cnt_l0_inc;
assign rsp_sft_cnt_l1_w = (layer_st) ? 8'h40   :
                          (dat_rsp_l1_stripe_end & ~dat_rsp_l1_block_end) ? rsp_sft_cnt_l1_ori :
                          (dat_rsp_l1_stripe_end & dat_rsp_l1_block_end) ? 8'h40   :
                          (dat_dummy_l1_en) ? (rsp_sft_cnt_l1_inc & 8'h3f) :
                          rsp_sft_cnt_l1_inc;
assign rsp_sft_cnt_l2_w = (layer_st) ? 8'h40   :
                          (dat_rsp_l2_stripe_end & ~dat_rsp_l2_block_end) ? rsp_sft_cnt_l2_ori :
                          (dat_rsp_l2_stripe_end & dat_rsp_l2_block_end) ? 8'h40   :
                          (dat_dummy_l2_en) ? (rsp_sft_cnt_l2_inc & 8'h3f) :
                          rsp_sft_cnt_l2_inc;
assign rsp_sft_cnt_l3_w = (layer_st) ? 8'h40   :
                          (dat_rsp_l3_stripe_end & ~dat_rsp_l3_block_end) ? rsp_sft_cnt_l3_ori :
                          (dat_rsp_l3_stripe_end & dat_rsp_l3_block_end) ? 8'h40   :
                          (dat_dummy_l3_en) ? (rsp_sft_cnt_l3_inc & 8'h3f) :
                          rsp_sft_cnt_l3_inc;
assign rsp_sft_cnt_l0_en = layer_st | (is_img_d1[17] & dat_rsp_l0_pvld);
assign rsp_sft_cnt_l1_en = layer_st | (is_img_d1[18] & dat_rsp_l1_pvld & (sub_h_total_g5 != 3'h1));
assign rsp_sft_cnt_l2_en = layer_st | (is_img_d1[19] & dat_rsp_l2_pvld & (sub_h_total_g5 == 3'h4));
assign rsp_sft_cnt_l3_en = layer_st | (is_img_d1[20] & dat_rsp_l3_pvld & (sub_h_total_g5 == 3'h4));
assign rsp_sft_cnt_l0_ori_en = layer_st | (is_img_d1[21] & dat_rsp_l0_pvld & dat_rsp_l0_stripe_end & dat_rsp_l0_block_end);
assign rsp_sft_cnt_l1_ori_en = layer_st | (is_img_d1[22] & dat_rsp_l1_pvld & dat_rsp_l1_stripe_end & dat_rsp_l1_block_end & (sub_h_total_g6 != 3'h1));
assign rsp_sft_cnt_l2_ori_en = layer_st | (is_img_d1[23] & dat_rsp_l2_pvld & dat_rsp_l2_stripe_end & dat_rsp_l2_block_end & (sub_h_total_g6 == 3'h4));
assign rsp_sft_cnt_l3_ori_en = layer_st | (is_img_d1[24] & dat_rsp_l3_pvld & dat_rsp_l3_stripe_end & dat_rsp_l3_block_end & (sub_h_total_g6 == 3'h4));
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l0_en\" -d \"rsp_sft_cnt_l0_w\" -q rsp_sft_cnt_l0");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l1_en\" -d \"rsp_sft_cnt_l1_w\" -q rsp_sft_cnt_l1");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l2_en\" -d \"rsp_sft_cnt_l2_w\" -q rsp_sft_cnt_l2");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l3_en\" -d \"rsp_sft_cnt_l3_w\" -q rsp_sft_cnt_l3");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l0_ori_en\" -d \"rsp_sft_cnt_l0_w\" -q rsp_sft_cnt_l0_ori");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l1_ori_en\" -d \"rsp_sft_cnt_l1_w\" -q rsp_sft_cnt_l1_ori");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l2_ori_en\" -d \"rsp_sft_cnt_l2_w\" -q rsp_sft_cnt_l2_ori");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l3_ori_en\" -d \"rsp_sft_cnt_l3_w\" -q rsp_sft_cnt_l3_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l0 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l0_en) == 1'b1) begin
           rsp_sft_cnt_l0 <= rsp_sft_cnt_l0_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l0_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l0 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l1 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l1_en) == 1'b1) begin
           rsp_sft_cnt_l1 <= rsp_sft_cnt_l1_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l1_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l2 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l2_en) == 1'b1) begin
           rsp_sft_cnt_l2 <= rsp_sft_cnt_l2_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l2_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l3 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l3_en) == 1'b1) begin
           rsp_sft_cnt_l3 <= rsp_sft_cnt_l3_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l3_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l0_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l0_ori_en) == 1'b1) begin
           rsp_sft_cnt_l0_ori <= rsp_sft_cnt_l0_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l0_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l0_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l1_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l1_ori_en) == 1'b1) begin
           rsp_sft_cnt_l1_ori <= rsp_sft_cnt_l1_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l1_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l1_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l2_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l2_ori_en) == 1'b1) begin
           rsp_sft_cnt_l2_ori <= rsp_sft_cnt_l2_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l2_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l2_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l3_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l3_ori_en) == 1'b1) begin
           rsp_sft_cnt_l3_ori <= rsp_sft_cnt_l3_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l3_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l3_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// response data                                      /////
//////////////////////////////////////////////////////////////
//////////////// data for winograd ////////////////
//winograd need future update

//////////////// data for convlution ////////////////
assign dat_rsp_pad_value = {64{pad_value[7:0]}};
assign dat_rsp_l0c0 = dat_l0c0_dummy ? dat_rsp_pad_value : dat_l0c0;
assign dat_rsp_l1c0 = dat_l1c0_dummy ? dat_rsp_pad_value : dat_l1c0;
assign dat_rsp_l2c0 = dat_l2c0_dummy ? dat_rsp_pad_value : dat_l2c0;
assign dat_rsp_l3c0 = dat_l3c0_dummy ? dat_rsp_pad_value : dat_l3c0;
assign dat_rsp_l0c1 = dat_l0c1_dummy ? dat_rsp_pad_value : dat_l0c1;
assign dat_rsp_l1c1 = dat_l1c1_dummy ? dat_rsp_pad_value : dat_l1c1;
assign dat_rsp_l2c1 = dat_l2c1_dummy ? dat_rsp_pad_value : dat_l2c1;
assign dat_rsp_l3c1 = dat_l3c1_dummy ? dat_rsp_pad_value : dat_l3c1;
//several atomM may combine together as an entry

assign dat_rsp_conv_8b = (is_winograd_d1[14] | is_img_d1[26]) ? {512{1'b0}} :
((dat_rsp_bytes <= 8'h20)&((dat_rsp_sub_w[0] == 1'h0))) ? {{512/2{1'b0}}, dat_rsp_l0c0[512/2 -1:0]} :
((dat_rsp_bytes <= 8'h20)&((dat_rsp_sub_w[0] == 1'h1))) ? {{512/2{1'b0}}, dat_rsp_l0c0[512 -1:512/2]} :
                dat_rsp_l0c0;
assign dat_rsp_conv = dat_rsp_conv_8b;
//////////////// data for image ////////////////
assign dat_rsp_l0_sft_in = ~is_img_d1[27] ? 'b0 : {dat_rsp_l0c0, dat_rsp_l0c1};
assign dat_rsp_l1_sft_in = ~is_img_d1[28] ? 'b0 : {dat_rsp_l1c0, dat_rsp_l1c1};
assign dat_rsp_l2_sft_in = ~is_img_d1[29] ? 'b0 : {dat_rsp_l2c0, dat_rsp_l2c1};
assign dat_rsp_l3_sft_in = ~is_img_d1[30] ? 'b0 : {dat_rsp_l3c0, dat_rsp_l3c1};
assign {mon_dat_rsp_l0_sft, dat_rsp_l0_sft} = dat_rsp_l0_sft_in >> {rsp_sft_cnt_l0, 3'b0};
assign {mon_dat_rsp_l1_sft, dat_rsp_l1_sft} = dat_rsp_l1_sft_in >> {rsp_sft_cnt_l1, 3'b0};
assign {mon_dat_rsp_l2_sft, dat_rsp_l2_sft} = dat_rsp_l2_sft_in >> {rsp_sft_cnt_l2, 3'b0};
assign {mon_dat_rsp_l3_sft, dat_rsp_l3_sft} = dat_rsp_l3_sft_in >> {rsp_sft_cnt_l3, 3'b0};
assign dat_rsp_img_8b = (~is_img_d1[32])? 'b0 :
                        (sub_h_total_g8 == 3'h4) ? {dat_rsp_l3_sft[512/4 -1:0], dat_rsp_l2_sft_d3[512/4 -1:0], dat_rsp_l1_sft_d3[512/4 -1:0], dat_rsp_l0_sft_d3[512/4 -1:0]} :
                        (sub_h_total_g8 == 3'h2) ? {dat_rsp_l1_sft[512/2 -1:0], dat_rsp_l0_sft_d1[512/2 -1:0]} :
                        dat_rsp_l0_sft[512 -1:0];
assign dat_rsp_img = dat_rsp_img_8b;
wire dat_rsp_sft_d1_en = dat_rsp_l0_pvld & (sub_h_total_g9 != 3'h1);
wire dat_rsp_sft_d2_en = dat_rsp_l1_pvld & (sub_h_total_g9 == 3'h4);
wire dat_rsp_sft_d3_en = dat_rsp_l2_pvld & (sub_h_total_g9 == 3'h4);
//: my $half=512/2;
//: my $quat=512/4;
//: &eperl::flop("-nodeclare -wid ${half} -norst -en \"dat_rsp_sft_d1_en\" -d \"dat_rsp_l0_sft\" -q dat_rsp_l0_sft_d1");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d2_en\" -d \"dat_rsp_l0_sft_d1\" -q dat_rsp_l0_sft_d2");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d3_en\" -d \"dat_rsp_l0_sft_d2\" -q dat_rsp_l0_sft_d3");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d2_en\" -d \"dat_rsp_l1_sft\" -q dat_rsp_l1_sft_d2");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d3_en\" -d \"dat_rsp_l1_sft_d2\" -q dat_rsp_l1_sft_d3");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d3_en\" -d \"dat_rsp_l2_sft\" -q dat_rsp_l2_sft_d3");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d1_en) == 1'b1) begin
           dat_rsp_l0_sft_d1 <= dat_rsp_l0_sft;
       // VCS coverage off
       end else if ((dat_rsp_sft_d1_en) == 1'b0) begin
       end else begin
           dat_rsp_l0_sft_d1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d2_en) == 1'b1) begin
           dat_rsp_l0_sft_d2 <= dat_rsp_l0_sft_d1;
       // VCS coverage off
       end else if ((dat_rsp_sft_d2_en) == 1'b0) begin
       end else begin
           dat_rsp_l0_sft_d2 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d3_en) == 1'b1) begin
           dat_rsp_l0_sft_d3 <= dat_rsp_l0_sft_d2;
       // VCS coverage off
       end else if ((dat_rsp_sft_d3_en) == 1'b0) begin
       end else begin
           dat_rsp_l0_sft_d3 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d2_en) == 1'b1) begin
           dat_rsp_l1_sft_d2 <= dat_rsp_l1_sft;
       // VCS coverage off
       end else if ((dat_rsp_sft_d2_en) == 1'b0) begin
       end else begin
           dat_rsp_l1_sft_d2 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d3_en) == 1'b1) begin
           dat_rsp_l1_sft_d3 <= dat_rsp_l1_sft_d2;
       // VCS coverage off
       end else if ((dat_rsp_sft_d3_en) == 1'b0) begin
       end else begin
           dat_rsp_l1_sft_d3 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d3_en) == 1'b1) begin
           dat_rsp_l2_sft_d3 <= dat_rsp_l2_sft;
       // VCS coverage off
       end else if ((dat_rsp_sft_d3_en) == 1'b0) begin
       end else begin
           dat_rsp_l2_sft_d3 <= 'bx;
       // VCS coverage on
       end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////// byte mask ////////////////
//sub_h_total=2, each sub_h align to 1/2 entry;
//sub_h_total=4, each sub_h align to 1/4 entry;
assign dat_rsp_ori_mask = ~({64{1'b1}} << dat_rsp_bytes);
assign dat_rsp_cur_h_mask_p1 = (dat_rsp_cur_sub_h >= 2'h1) ? {64{1'b1}} : 'b0;
assign dat_rsp_cur_h_mask_p2 = (dat_rsp_cur_sub_h >= 2'h2) ? {64/2{1'b1}} : 'b0;
assign dat_rsp_cur_h_mask_p3 = (dat_rsp_cur_sub_h == 2'h3) ? {64/2{1'b1}} : 'b0;
assign dat_rsp_cur_h_e2_mask_8b = {dat_rsp_cur_h_mask_p1[64/2 -1:0], {64/2{1'b1}}};
assign dat_rsp_cur_h_e4_mask_8b = {dat_rsp_cur_h_mask_p3[64/4 -1:0], dat_rsp_cur_h_mask_p2[64/4 -1:0], dat_rsp_cur_h_mask_p1[64/4 -1:0], {64/4{1'b1}}};
assign dat_rsp_mask_8b = (sub_h_total_g11 == 3'h4) ? ({4{dat_rsp_ori_mask[64/4 -1:0]}} & dat_rsp_cur_h_e4_mask_8b) :
                         (sub_h_total_g11 == 3'h2) ? ({2{dat_rsp_ori_mask[64/2 -1:0]}} & dat_rsp_cur_h_e2_mask_8b) :
                         dat_rsp_ori_mask[64 -1:0];
assign dat_rsp_data_w = is_img_d1[33] ? dat_rsp_img :
                        dat_rsp_conv;
//: my $i;
//: my $b1;
//: my $b0;
//: my $kk=64 -1;
//: print "assign dat_rsp_mask_val_int8 = {";
//: for($i = ${kk}; $i >= 0; $i --) {
//: $b0 = sprintf("%3d", $i * 8);
//: $b1 = sprintf("%3d", $i * 8 + 7);
//: print "(|dat_rsp_data_w[${b1}:${b0}])";
//: if($i == 0) {
//: print "};\n";
//: } elsif ($i % 8 == 0) {
//: print ",\n                               ";
//: } else {
//: print ", ";
//: }
//: }
//: print "\n\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_rsp_mask_val_int8 = {(|dat_rsp_data_w[511:504]), (|dat_rsp_data_w[503:496]), (|dat_rsp_data_w[495:488]), (|dat_rsp_data_w[487:480]), (|dat_rsp_data_w[479:472]), (|dat_rsp_data_w[471:464]), (|dat_rsp_data_w[463:456]), (|dat_rsp_data_w[455:448]),
                               (|dat_rsp_data_w[447:440]), (|dat_rsp_data_w[439:432]), (|dat_rsp_data_w[431:424]), (|dat_rsp_data_w[423:416]), (|dat_rsp_data_w[415:408]), (|dat_rsp_data_w[407:400]), (|dat_rsp_data_w[399:392]), (|dat_rsp_data_w[391:384]),
                               (|dat_rsp_data_w[383:376]), (|dat_rsp_data_w[375:368]), (|dat_rsp_data_w[367:360]), (|dat_rsp_data_w[359:352]), (|dat_rsp_data_w[351:344]), (|dat_rsp_data_w[343:336]), (|dat_rsp_data_w[335:328]), (|dat_rsp_data_w[327:320]),
                               (|dat_rsp_data_w[319:312]), (|dat_rsp_data_w[311:304]), (|dat_rsp_data_w[303:296]), (|dat_rsp_data_w[295:288]), (|dat_rsp_data_w[287:280]), (|dat_rsp_data_w[279:272]), (|dat_rsp_data_w[271:264]), (|dat_rsp_data_w[263:256]),
                               (|dat_rsp_data_w[255:248]), (|dat_rsp_data_w[247:240]), (|dat_rsp_data_w[239:232]), (|dat_rsp_data_w[231:224]), (|dat_rsp_data_w[223:216]), (|dat_rsp_data_w[215:208]), (|dat_rsp_data_w[207:200]), (|dat_rsp_data_w[199:192]),
                               (|dat_rsp_data_w[191:184]), (|dat_rsp_data_w[183:176]), (|dat_rsp_data_w[175:168]), (|dat_rsp_data_w[167:160]), (|dat_rsp_data_w[159:152]), (|dat_rsp_data_w[151:144]), (|dat_rsp_data_w[143:136]), (|dat_rsp_data_w[135:128]),
                               (|dat_rsp_data_w[127:120]), (|dat_rsp_data_w[119:112]), (|dat_rsp_data_w[111:104]), (|dat_rsp_data_w[103: 96]), (|dat_rsp_data_w[ 95: 88]), (|dat_rsp_data_w[ 87: 80]), (|dat_rsp_data_w[ 79: 72]), (|dat_rsp_data_w[ 71: 64]),
                               (|dat_rsp_data_w[ 63: 56]), (|dat_rsp_data_w[ 55: 48]), (|dat_rsp_data_w[ 47: 40]), (|dat_rsp_data_w[ 39: 32]), (|dat_rsp_data_w[ 31: 24]), (|dat_rsp_data_w[ 23: 16]), (|dat_rsp_data_w[ 15:  8]), (|dat_rsp_data_w[  7:  0])};



//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dat_rsp_mask_w = (dat_rsp_mask_8b & dat_rsp_mask_val_int8) ;
assign dat_rsp_p1_vld_w = 1'b0;
assign dat_rsp_p0_vld_w = dat_rsp_pvld & ~is_winograd_d1[16];
//////////////////////////////////////////////////////////////
///// latency register to balance with PRA cell          /////
//////////////////////////////////////////////////////////////
//: my $total_latency = 5;
//:
//: print "assign dat_out_pvld_l0 = dat_rsp_pvld;\n";
//: print "assign dat_out_flag_l0 = dat_rsp_flag;\n";
//: for(my $i = 0; $i < $total_latency; $i ++) {
//: my $j = $i + 1;
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -d \"dat_out_pvld_l${i}\"   -q dat_out_pvld_l${j}");
//: &eperl::flop("-wid 9   -rval \"{9{1'b0}}\"  -en \"dat_out_pvld_l${i}\"  -d \"dat_out_flag_l${i}\" -q dat_out_flag_l${j}");
//: }
//:
//: my $k = $total_latency;
//: print "assign dat_out_pvld_w = is_winograd_d1[17] ? dat_out_pvld_l${k} : dat_rsp_pvld;\n";
//: print "assign dat_out_flag_w = is_winograd_d1[18] ? dat_out_flag_l${k} : dat_rsp_flag;\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_out_pvld_l0 = dat_rsp_pvld;
assign dat_out_flag_l0 = dat_rsp_flag;
reg  dat_out_pvld_l1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l1 <= 1'b0;
   end else begin
       dat_out_pvld_l1 <= dat_out_pvld_l0;
   end
end
reg [8:0] dat_out_flag_l1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l1 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l0) == 1'b1) begin
           dat_out_flag_l1 <= dat_out_flag_l0;
       // VCS coverage off
       end else if ((dat_out_pvld_l0) == 1'b0) begin
       end else begin
           dat_out_flag_l1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l2 <= 1'b0;
   end else begin
       dat_out_pvld_l2 <= dat_out_pvld_l1;
   end
end
reg [8:0] dat_out_flag_l2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l2 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l1) == 1'b1) begin
           dat_out_flag_l2 <= dat_out_flag_l1;
       // VCS coverage off
       end else if ((dat_out_pvld_l1) == 1'b0) begin
       end else begin
           dat_out_flag_l2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l3 <= 1'b0;
   end else begin
       dat_out_pvld_l3 <= dat_out_pvld_l2;
   end
end
reg [8:0] dat_out_flag_l3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l3 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l2) == 1'b1) begin
           dat_out_flag_l3 <= dat_out_flag_l2;
       // VCS coverage off
       end else if ((dat_out_pvld_l2) == 1'b0) begin
       end else begin
           dat_out_flag_l3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l4 <= 1'b0;
   end else begin
       dat_out_pvld_l4 <= dat_out_pvld_l3;
   end
end
reg [8:0] dat_out_flag_l4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l4 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l3) == 1'b1) begin
           dat_out_flag_l4 <= dat_out_flag_l3;
       // VCS coverage off
       end else if ((dat_out_pvld_l3) == 1'b0) begin
       end else begin
           dat_out_flag_l4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l5 <= 1'b0;
   end else begin
       dat_out_pvld_l5 <= dat_out_pvld_l4;
   end
end
reg [8:0] dat_out_flag_l5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l5 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l4) == 1'b1) begin
           dat_out_flag_l5 <= dat_out_flag_l4;
       // VCS coverage off
       end else if ((dat_out_pvld_l4) == 1'b0) begin
       end else begin
           dat_out_flag_l5 <= 'bx;
       // VCS coverage on
       end
   end
end
assign dat_out_pvld_w = is_winograd_d1[17] ? dat_out_pvld_l5 : dat_rsp_pvld;
assign dat_out_flag_w = is_winograd_d1[18] ? dat_out_flag_l5 : dat_rsp_flag;

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dat_out_bypass_p0_vld_w = dat_rsp_p0_vld_w;
assign dat_out_bypass_mask_w = dat_rsp_mask_w;
assign dat_out_bypass_data_w = dat_rsp_data_w;
//: my $kk=64;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_out_pvld_w\" -q dat_out_pvld");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_out_pvld_w\" -d \"dat_out_flag_w\" -q dat_out_flag");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dat_out_bypass_p0_vld_w\" -d \"dat_out_bypass_mask_w\" -q dat_out_bypass_mask");
//: for(my $i = 0; $i < 64; $i ++) {
//: my $b0 = $i * 8;
//: my $b1 = $i * 8 + 7;
//: &eperl::flop("-nodeclare  -norst -en \"dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[${i}]\" -d \"dat_out_bypass_data_w[${b1}:${b0}]\" -q dat_out_bypass_data[${b1}:${b0}]");
//: }
//:
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld <= 1'b0;
   end else begin
       dat_out_pvld <= dat_out_pvld_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_w) == 1'b1) begin
           dat_out_flag <= dat_out_flag_w;
       // VCS coverage off
       end else if ((dat_out_pvld_w) == 1'b0) begin
       end else begin
           dat_out_flag <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_bypass_mask <= {64{1'b0}};
   end else begin
       if ((dat_out_bypass_p0_vld_w) == 1'b1) begin
           dat_out_bypass_mask <= dat_out_bypass_mask_w;
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w) == 1'b0) begin
       end else begin
           dat_out_bypass_mask <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[0]) == 1'b1) begin
           dat_out_bypass_data[7:0] <= dat_out_bypass_data_w[7:0];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[0]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[7:0] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[1]) == 1'b1) begin
           dat_out_bypass_data[15:8] <= dat_out_bypass_data_w[15:8];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[1]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[15:8] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[2]) == 1'b1) begin
           dat_out_bypass_data[23:16] <= dat_out_bypass_data_w[23:16];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[2]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[23:16] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[3]) == 1'b1) begin
           dat_out_bypass_data[31:24] <= dat_out_bypass_data_w[31:24];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[3]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[31:24] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[4]) == 1'b1) begin
           dat_out_bypass_data[39:32] <= dat_out_bypass_data_w[39:32];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[4]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[39:32] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[5]) == 1'b1) begin
           dat_out_bypass_data[47:40] <= dat_out_bypass_data_w[47:40];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[5]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[47:40] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[6]) == 1'b1) begin
           dat_out_bypass_data[55:48] <= dat_out_bypass_data_w[55:48];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[6]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[55:48] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[7]) == 1'b1) begin
           dat_out_bypass_data[63:56] <= dat_out_bypass_data_w[63:56];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[7]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[63:56] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[8]) == 1'b1) begin
           dat_out_bypass_data[71:64] <= dat_out_bypass_data_w[71:64];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[8]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[71:64] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[9]) == 1'b1) begin
           dat_out_bypass_data[79:72] <= dat_out_bypass_data_w[79:72];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[9]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[79:72] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[10]) == 1'b1) begin
           dat_out_bypass_data[87:80] <= dat_out_bypass_data_w[87:80];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[10]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[87:80] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[11]) == 1'b1) begin
           dat_out_bypass_data[95:88] <= dat_out_bypass_data_w[95:88];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[11]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[95:88] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[12]) == 1'b1) begin
           dat_out_bypass_data[103:96] <= dat_out_bypass_data_w[103:96];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[12]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[103:96] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[13]) == 1'b1) begin
           dat_out_bypass_data[111:104] <= dat_out_bypass_data_w[111:104];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[13]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[111:104] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[14]) == 1'b1) begin
           dat_out_bypass_data[119:112] <= dat_out_bypass_data_w[119:112];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[14]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[119:112] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[15]) == 1'b1) begin
           dat_out_bypass_data[127:120] <= dat_out_bypass_data_w[127:120];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[15]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[127:120] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[16]) == 1'b1) begin
           dat_out_bypass_data[135:128] <= dat_out_bypass_data_w[135:128];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[16]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[135:128] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[17]) == 1'b1) begin
           dat_out_bypass_data[143:136] <= dat_out_bypass_data_w[143:136];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[17]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[143:136] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[18]) == 1'b1) begin
           dat_out_bypass_data[151:144] <= dat_out_bypass_data_w[151:144];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[18]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[151:144] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[19]) == 1'b1) begin
           dat_out_bypass_data[159:152] <= dat_out_bypass_data_w[159:152];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[19]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[159:152] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[20]) == 1'b1) begin
           dat_out_bypass_data[167:160] <= dat_out_bypass_data_w[167:160];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[20]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[167:160] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[21]) == 1'b1) begin
           dat_out_bypass_data[175:168] <= dat_out_bypass_data_w[175:168];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[21]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[175:168] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[22]) == 1'b1) begin
           dat_out_bypass_data[183:176] <= dat_out_bypass_data_w[183:176];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[22]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[183:176] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[23]) == 1'b1) begin
           dat_out_bypass_data[191:184] <= dat_out_bypass_data_w[191:184];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[23]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[191:184] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[24]) == 1'b1) begin
           dat_out_bypass_data[199:192] <= dat_out_bypass_data_w[199:192];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[24]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[199:192] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[25]) == 1'b1) begin
           dat_out_bypass_data[207:200] <= dat_out_bypass_data_w[207:200];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[25]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[207:200] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[26]) == 1'b1) begin
           dat_out_bypass_data[215:208] <= dat_out_bypass_data_w[215:208];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[26]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[215:208] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[27]) == 1'b1) begin
           dat_out_bypass_data[223:216] <= dat_out_bypass_data_w[223:216];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[27]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[223:216] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[28]) == 1'b1) begin
           dat_out_bypass_data[231:224] <= dat_out_bypass_data_w[231:224];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[28]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[231:224] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[29]) == 1'b1) begin
           dat_out_bypass_data[239:232] <= dat_out_bypass_data_w[239:232];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[29]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[239:232] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[30]) == 1'b1) begin
           dat_out_bypass_data[247:240] <= dat_out_bypass_data_w[247:240];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[30]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[247:240] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[31]) == 1'b1) begin
           dat_out_bypass_data[255:248] <= dat_out_bypass_data_w[255:248];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[31]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[255:248] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[32]) == 1'b1) begin
           dat_out_bypass_data[263:256] <= dat_out_bypass_data_w[263:256];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[32]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[263:256] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[33]) == 1'b1) begin
           dat_out_bypass_data[271:264] <= dat_out_bypass_data_w[271:264];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[33]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[271:264] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[34]) == 1'b1) begin
           dat_out_bypass_data[279:272] <= dat_out_bypass_data_w[279:272];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[34]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[279:272] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[35]) == 1'b1) begin
           dat_out_bypass_data[287:280] <= dat_out_bypass_data_w[287:280];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[35]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[287:280] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[36]) == 1'b1) begin
           dat_out_bypass_data[295:288] <= dat_out_bypass_data_w[295:288];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[36]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[295:288] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[37]) == 1'b1) begin
           dat_out_bypass_data[303:296] <= dat_out_bypass_data_w[303:296];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[37]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[303:296] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[38]) == 1'b1) begin
           dat_out_bypass_data[311:304] <= dat_out_bypass_data_w[311:304];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[38]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[311:304] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[39]) == 1'b1) begin
           dat_out_bypass_data[319:312] <= dat_out_bypass_data_w[319:312];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[39]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[319:312] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[40]) == 1'b1) begin
           dat_out_bypass_data[327:320] <= dat_out_bypass_data_w[327:320];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[40]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[327:320] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[41]) == 1'b1) begin
           dat_out_bypass_data[335:328] <= dat_out_bypass_data_w[335:328];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[41]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[335:328] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[42]) == 1'b1) begin
           dat_out_bypass_data[343:336] <= dat_out_bypass_data_w[343:336];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[42]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[343:336] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[43]) == 1'b1) begin
           dat_out_bypass_data[351:344] <= dat_out_bypass_data_w[351:344];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[43]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[351:344] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[44]) == 1'b1) begin
           dat_out_bypass_data[359:352] <= dat_out_bypass_data_w[359:352];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[44]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[359:352] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[45]) == 1'b1) begin
           dat_out_bypass_data[367:360] <= dat_out_bypass_data_w[367:360];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[45]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[367:360] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[46]) == 1'b1) begin
           dat_out_bypass_data[375:368] <= dat_out_bypass_data_w[375:368];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[46]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[375:368] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[47]) == 1'b1) begin
           dat_out_bypass_data[383:376] <= dat_out_bypass_data_w[383:376];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[47]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[383:376] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[48]) == 1'b1) begin
           dat_out_bypass_data[391:384] <= dat_out_bypass_data_w[391:384];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[48]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[391:384] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[49]) == 1'b1) begin
           dat_out_bypass_data[399:392] <= dat_out_bypass_data_w[399:392];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[49]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[399:392] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[50]) == 1'b1) begin
           dat_out_bypass_data[407:400] <= dat_out_bypass_data_w[407:400];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[50]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[407:400] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[51]) == 1'b1) begin
           dat_out_bypass_data[415:408] <= dat_out_bypass_data_w[415:408];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[51]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[415:408] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[52]) == 1'b1) begin
           dat_out_bypass_data[423:416] <= dat_out_bypass_data_w[423:416];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[52]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[423:416] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[53]) == 1'b1) begin
           dat_out_bypass_data[431:424] <= dat_out_bypass_data_w[431:424];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[53]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[431:424] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[54]) == 1'b1) begin
           dat_out_bypass_data[439:432] <= dat_out_bypass_data_w[439:432];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[54]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[439:432] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[55]) == 1'b1) begin
           dat_out_bypass_data[447:440] <= dat_out_bypass_data_w[447:440];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[55]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[447:440] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[56]) == 1'b1) begin
           dat_out_bypass_data[455:448] <= dat_out_bypass_data_w[455:448];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[56]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[455:448] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[57]) == 1'b1) begin
           dat_out_bypass_data[463:456] <= dat_out_bypass_data_w[463:456];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[57]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[463:456] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[58]) == 1'b1) begin
           dat_out_bypass_data[471:464] <= dat_out_bypass_data_w[471:464];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[58]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[471:464] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[59]) == 1'b1) begin
           dat_out_bypass_data[479:472] <= dat_out_bypass_data_w[479:472];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[59]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[479:472] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[60]) == 1'b1) begin
           dat_out_bypass_data[487:480] <= dat_out_bypass_data_w[487:480];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[60]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[487:480] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[61]) == 1'b1) begin
           dat_out_bypass_data[495:488] <= dat_out_bypass_data_w[495:488];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[61]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[495:488] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[62]) == 1'b1) begin
           dat_out_bypass_data[503:496] <= dat_out_bypass_data_w[503:496];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[62]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[503:496] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[63]) == 1'b1) begin
           dat_out_bypass_data[511:504] <= dat_out_bypass_data_w[511:504];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[63]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[511:504] <= 'bx;
       // VCS coverage on
       end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)

assign dat_out_wg_data = {512{1'b0}};
assign dat_out_wg_mask = {64{1'b0}};
//////////////////////////////////////////////////////////////
///// finial registers                                   /////
//////////////////////////////////////////////////////////////
assign dat_out_data = is_winograd_d1[20] ? dat_out_wg_data : dat_out_bypass_data;
assign dat_out_mask = ~dat_out_pvld ? 'b0 : is_winograd_d1[21] ? dat_out_wg_mask : dat_out_bypass_mask;
//: my $kk=64;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_out_pvld\" -q dl_out_pvld");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dat_out_pvld | dl_out_pvld\" -d \"dat_out_mask\" -q dl_out_mask");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_out_pvld\" -d \"dat_out_flag\" -q dl_out_flag");
//: my $i;
//: my $b0;
//: my $b1;
//: my $kk= 8;
//: for($i = 0; $i < 64; $i ++) {
//: $b0 = $i * 8;
//: $b1 = $i * 8 + 7;
//: &eperl::flop("-wid ${kk}  -norst -en \"dat_out_mask[$i]\" -d \"dat_out_data[${b1}:${b0}]\" -q dl_out_data${i}");
//: }
//: print "\n\n\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_pvld <= 1'b0;
   end else begin
       dl_out_pvld <= dat_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_mask <= {64{1'b0}};
   end else begin
       if ((dat_out_pvld | dl_out_pvld) == 1'b1) begin
           dl_out_mask <= dat_out_mask;
       // VCS coverage off
       end else if ((dat_out_pvld | dl_out_pvld) == 1'b0) begin
       end else begin
           dl_out_mask <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_flag <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld) == 1'b1) begin
           dl_out_flag <= dat_out_flag;
       // VCS coverage off
       end else if ((dat_out_pvld) == 1'b0) begin
       end else begin
           dl_out_flag <= 'bx;
       // VCS coverage on
       end
   end
end
reg [7:0] dl_out_data0;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[0]) == 1'b1) begin
           dl_out_data0 <= dat_out_data[7:0];
       // VCS coverage off
       end else if ((dat_out_mask[0]) == 1'b0) begin
       end else begin
           dl_out_data0 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data1;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[1]) == 1'b1) begin
           dl_out_data1 <= dat_out_data[15:8];
       // VCS coverage off
       end else if ((dat_out_mask[1]) == 1'b0) begin
       end else begin
           dl_out_data1 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data2;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[2]) == 1'b1) begin
           dl_out_data2 <= dat_out_data[23:16];
       // VCS coverage off
       end else if ((dat_out_mask[2]) == 1'b0) begin
       end else begin
           dl_out_data2 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data3;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[3]) == 1'b1) begin
           dl_out_data3 <= dat_out_data[31:24];
       // VCS coverage off
       end else if ((dat_out_mask[3]) == 1'b0) begin
       end else begin
           dl_out_data3 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data4;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[4]) == 1'b1) begin
           dl_out_data4 <= dat_out_data[39:32];
       // VCS coverage off
       end else if ((dat_out_mask[4]) == 1'b0) begin
       end else begin
           dl_out_data4 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data5;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[5]) == 1'b1) begin
           dl_out_data5 <= dat_out_data[47:40];
       // VCS coverage off
       end else if ((dat_out_mask[5]) == 1'b0) begin
       end else begin
           dl_out_data5 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data6;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[6]) == 1'b1) begin
           dl_out_data6 <= dat_out_data[55:48];
       // VCS coverage off
       end else if ((dat_out_mask[6]) == 1'b0) begin
       end else begin
           dl_out_data6 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data7;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[7]) == 1'b1) begin
           dl_out_data7 <= dat_out_data[63:56];
       // VCS coverage off
       end else if ((dat_out_mask[7]) == 1'b0) begin
       end else begin
           dl_out_data7 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data8;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[8]) == 1'b1) begin
           dl_out_data8 <= dat_out_data[71:64];
       // VCS coverage off
       end else if ((dat_out_mask[8]) == 1'b0) begin
       end else begin
           dl_out_data8 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data9;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[9]) == 1'b1) begin
           dl_out_data9 <= dat_out_data[79:72];
       // VCS coverage off
       end else if ((dat_out_mask[9]) == 1'b0) begin
       end else begin
           dl_out_data9 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data10;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[10]) == 1'b1) begin
           dl_out_data10 <= dat_out_data[87:80];
       // VCS coverage off
       end else if ((dat_out_mask[10]) == 1'b0) begin
       end else begin
           dl_out_data10 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data11;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[11]) == 1'b1) begin
           dl_out_data11 <= dat_out_data[95:88];
       // VCS coverage off
       end else if ((dat_out_mask[11]) == 1'b0) begin
       end else begin
           dl_out_data11 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data12;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[12]) == 1'b1) begin
           dl_out_data12 <= dat_out_data[103:96];
       // VCS coverage off
       end else if ((dat_out_mask[12]) == 1'b0) begin
       end else begin
           dl_out_data12 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data13;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[13]) == 1'b1) begin
           dl_out_data13 <= dat_out_data[111:104];
       // VCS coverage off
       end else if ((dat_out_mask[13]) == 1'b0) begin
       end else begin
           dl_out_data13 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data14;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[14]) == 1'b1) begin
           dl_out_data14 <= dat_out_data[119:112];
       // VCS coverage off
       end else if ((dat_out_mask[14]) == 1'b0) begin
       end else begin
           dl_out_data14 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data15;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[15]) == 1'b1) begin
           dl_out_data15 <= dat_out_data[127:120];
       // VCS coverage off
       end else if ((dat_out_mask[15]) == 1'b0) begin
       end else begin
           dl_out_data15 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data16;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[16]) == 1'b1) begin
           dl_out_data16 <= dat_out_data[135:128];
       // VCS coverage off
       end else if ((dat_out_mask[16]) == 1'b0) begin
       end else begin
           dl_out_data16 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data17;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[17]) == 1'b1) begin
           dl_out_data17 <= dat_out_data[143:136];
       // VCS coverage off
       end else if ((dat_out_mask[17]) == 1'b0) begin
       end else begin
           dl_out_data17 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data18;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[18]) == 1'b1) begin
           dl_out_data18 <= dat_out_data[151:144];
       // VCS coverage off
       end else if ((dat_out_mask[18]) == 1'b0) begin
       end else begin
           dl_out_data18 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data19;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[19]) == 1'b1) begin
           dl_out_data19 <= dat_out_data[159:152];
       // VCS coverage off
       end else if ((dat_out_mask[19]) == 1'b0) begin
       end else begin
           dl_out_data19 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data20;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[20]) == 1'b1) begin
           dl_out_data20 <= dat_out_data[167:160];
       // VCS coverage off
       end else if ((dat_out_mask[20]) == 1'b0) begin
       end else begin
           dl_out_data20 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data21;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[21]) == 1'b1) begin
           dl_out_data21 <= dat_out_data[175:168];
       // VCS coverage off
       end else if ((dat_out_mask[21]) == 1'b0) begin
       end else begin
           dl_out_data21 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data22;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[22]) == 1'b1) begin
           dl_out_data22 <= dat_out_data[183:176];
       // VCS coverage off
       end else if ((dat_out_mask[22]) == 1'b0) begin
       end else begin
           dl_out_data22 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data23;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[23]) == 1'b1) begin
           dl_out_data23 <= dat_out_data[191:184];
       // VCS coverage off
       end else if ((dat_out_mask[23]) == 1'b0) begin
       end else begin
           dl_out_data23 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data24;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[24]) == 1'b1) begin
           dl_out_data24 <= dat_out_data[199:192];
       // VCS coverage off
       end else if ((dat_out_mask[24]) == 1'b0) begin
       end else begin
           dl_out_data24 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data25;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[25]) == 1'b1) begin
           dl_out_data25 <= dat_out_data[207:200];
       // VCS coverage off
       end else if ((dat_out_mask[25]) == 1'b0) begin
       end else begin
           dl_out_data25 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data26;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[26]) == 1'b1) begin
           dl_out_data26 <= dat_out_data[215:208];
       // VCS coverage off
       end else if ((dat_out_mask[26]) == 1'b0) begin
       end else begin
           dl_out_data26 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data27;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[27]) == 1'b1) begin
           dl_out_data27 <= dat_out_data[223:216];
       // VCS coverage off
       end else if ((dat_out_mask[27]) == 1'b0) begin
       end else begin
           dl_out_data27 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data28;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[28]) == 1'b1) begin
           dl_out_data28 <= dat_out_data[231:224];
       // VCS coverage off
       end else if ((dat_out_mask[28]) == 1'b0) begin
       end else begin
           dl_out_data28 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data29;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[29]) == 1'b1) begin
           dl_out_data29 <= dat_out_data[239:232];
       // VCS coverage off
       end else if ((dat_out_mask[29]) == 1'b0) begin
       end else begin
           dl_out_data29 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data30;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[30]) == 1'b1) begin
           dl_out_data30 <= dat_out_data[247:240];
       // VCS coverage off
       end else if ((dat_out_mask[30]) == 1'b0) begin
       end else begin
           dl_out_data30 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data31;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[31]) == 1'b1) begin
           dl_out_data31 <= dat_out_data[255:248];
       // VCS coverage off
       end else if ((dat_out_mask[31]) == 1'b0) begin
       end else begin
           dl_out_data31 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data32;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[32]) == 1'b1) begin
           dl_out_data32 <= dat_out_data[263:256];
       // VCS coverage off
       end else if ((dat_out_mask[32]) == 1'b0) begin
       end else begin
           dl_out_data32 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data33;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[33]) == 1'b1) begin
           dl_out_data33 <= dat_out_data[271:264];
       // VCS coverage off
       end else if ((dat_out_mask[33]) == 1'b0) begin
       end else begin
           dl_out_data33 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data34;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[34]) == 1'b1) begin
           dl_out_data34 <= dat_out_data[279:272];
       // VCS coverage off
       end else if ((dat_out_mask[34]) == 1'b0) begin
       end else begin
           dl_out_data34 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data35;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[35]) == 1'b1) begin
           dl_out_data35 <= dat_out_data[287:280];
       // VCS coverage off
       end else if ((dat_out_mask[35]) == 1'b0) begin
       end else begin
           dl_out_data35 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data36;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[36]) == 1'b1) begin
           dl_out_data36 <= dat_out_data[295:288];
       // VCS coverage off
       end else if ((dat_out_mask[36]) == 1'b0) begin
       end else begin
           dl_out_data36 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data37;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[37]) == 1'b1) begin
           dl_out_data37 <= dat_out_data[303:296];
       // VCS coverage off
       end else if ((dat_out_mask[37]) == 1'b0) begin
       end else begin
           dl_out_data37 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data38;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[38]) == 1'b1) begin
           dl_out_data38 <= dat_out_data[311:304];
       // VCS coverage off
       end else if ((dat_out_mask[38]) == 1'b0) begin
       end else begin
           dl_out_data38 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data39;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[39]) == 1'b1) begin
           dl_out_data39 <= dat_out_data[319:312];
       // VCS coverage off
       end else if ((dat_out_mask[39]) == 1'b0) begin
       end else begin
           dl_out_data39 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data40;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[40]) == 1'b1) begin
           dl_out_data40 <= dat_out_data[327:320];
       // VCS coverage off
       end else if ((dat_out_mask[40]) == 1'b0) begin
       end else begin
           dl_out_data40 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data41;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[41]) == 1'b1) begin
           dl_out_data41 <= dat_out_data[335:328];
       // VCS coverage off
       end else if ((dat_out_mask[41]) == 1'b0) begin
       end else begin
           dl_out_data41 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data42;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[42]) == 1'b1) begin
           dl_out_data42 <= dat_out_data[343:336];
       // VCS coverage off
       end else if ((dat_out_mask[42]) == 1'b0) begin
       end else begin
           dl_out_data42 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data43;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[43]) == 1'b1) begin
           dl_out_data43 <= dat_out_data[351:344];
       // VCS coverage off
       end else if ((dat_out_mask[43]) == 1'b0) begin
       end else begin
           dl_out_data43 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data44;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[44]) == 1'b1) begin
           dl_out_data44 <= dat_out_data[359:352];
       // VCS coverage off
       end else if ((dat_out_mask[44]) == 1'b0) begin
       end else begin
           dl_out_data44 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data45;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[45]) == 1'b1) begin
           dl_out_data45 <= dat_out_data[367:360];
       // VCS coverage off
       end else if ((dat_out_mask[45]) == 1'b0) begin
       end else begin
           dl_out_data45 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data46;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[46]) == 1'b1) begin
           dl_out_data46 <= dat_out_data[375:368];
       // VCS coverage off
       end else if ((dat_out_mask[46]) == 1'b0) begin
       end else begin
           dl_out_data46 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data47;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[47]) == 1'b1) begin
           dl_out_data47 <= dat_out_data[383:376];
       // VCS coverage off
       end else if ((dat_out_mask[47]) == 1'b0) begin
       end else begin
           dl_out_data47 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data48;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[48]) == 1'b1) begin
           dl_out_data48 <= dat_out_data[391:384];
       // VCS coverage off
       end else if ((dat_out_mask[48]) == 1'b0) begin
       end else begin
           dl_out_data48 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data49;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[49]) == 1'b1) begin
           dl_out_data49 <= dat_out_data[399:392];
       // VCS coverage off
       end else if ((dat_out_mask[49]) == 1'b0) begin
       end else begin
           dl_out_data49 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data50;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[50]) == 1'b1) begin
           dl_out_data50 <= dat_out_data[407:400];
       // VCS coverage off
       end else if ((dat_out_mask[50]) == 1'b0) begin
       end else begin
           dl_out_data50 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data51;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[51]) == 1'b1) begin
           dl_out_data51 <= dat_out_data[415:408];
       // VCS coverage off
       end else if ((dat_out_mask[51]) == 1'b0) begin
       end else begin
           dl_out_data51 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data52;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[52]) == 1'b1) begin
           dl_out_data52 <= dat_out_data[423:416];
       // VCS coverage off
       end else if ((dat_out_mask[52]) == 1'b0) begin
       end else begin
           dl_out_data52 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data53;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[53]) == 1'b1) begin
           dl_out_data53 <= dat_out_data[431:424];
       // VCS coverage off
       end else if ((dat_out_mask[53]) == 1'b0) begin
       end else begin
           dl_out_data53 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data54;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[54]) == 1'b1) begin
           dl_out_data54 <= dat_out_data[439:432];
       // VCS coverage off
       end else if ((dat_out_mask[54]) == 1'b0) begin
       end else begin
           dl_out_data54 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data55;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[55]) == 1'b1) begin
           dl_out_data55 <= dat_out_data[447:440];
       // VCS coverage off
       end else if ((dat_out_mask[55]) == 1'b0) begin
       end else begin
           dl_out_data55 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data56;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[56]) == 1'b1) begin
           dl_out_data56 <= dat_out_data[455:448];
       // VCS coverage off
       end else if ((dat_out_mask[56]) == 1'b0) begin
       end else begin
           dl_out_data56 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data57;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[57]) == 1'b1) begin
           dl_out_data57 <= dat_out_data[463:456];
       // VCS coverage off
       end else if ((dat_out_mask[57]) == 1'b0) begin
       end else begin
           dl_out_data57 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data58;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[58]) == 1'b1) begin
           dl_out_data58 <= dat_out_data[471:464];
       // VCS coverage off
       end else if ((dat_out_mask[58]) == 1'b0) begin
       end else begin
           dl_out_data58 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data59;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[59]) == 1'b1) begin
           dl_out_data59 <= dat_out_data[479:472];
       // VCS coverage off
       end else if ((dat_out_mask[59]) == 1'b0) begin
       end else begin
           dl_out_data59 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data60;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[60]) == 1'b1) begin
           dl_out_data60 <= dat_out_data[487:480];
       // VCS coverage off
       end else if ((dat_out_mask[60]) == 1'b0) begin
       end else begin
           dl_out_data60 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data61;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[61]) == 1'b1) begin
           dl_out_data61 <= dat_out_data[495:488];
       // VCS coverage off
       end else if ((dat_out_mask[61]) == 1'b0) begin
       end else begin
           dl_out_data61 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data62;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[62]) == 1'b1) begin
           dl_out_data62 <= dat_out_data[503:496];
       // VCS coverage off
       end else if ((dat_out_mask[62]) == 1'b0) begin
       end else begin
           dl_out_data62 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data63;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[63]) == 1'b1) begin
           dl_out_data63 <= dat_out_data[511:504];
       // VCS coverage off
       end else if ((dat_out_mask[63]) == 1'b0) begin
       end else begin
           dl_out_data63 <= 'bx;
       // VCS coverage on
       end
end




//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// registers for retiming                             /////
//////////////////////////////////////////////////////////////
assign sc2mac_dat_pd_w = ~dl_out_pvld ? 9'b0 : dl_out_flag;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dl_out_pvld\" -q dl_out_pvld_d1");
//: my $kk=64;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dl_out_pvld\" -q sc2mac_dat_a_pvld");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dl_out_pvld\" -q sc2mac_dat_b_pvld");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"sc2mac_dat_pd_w\" -q sc2mac_dat_a_pd");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"sc2mac_dat_pd_w\" -q sc2mac_dat_b_pd");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"dl_out_mask\" -q sc2mac_dat_a_mask");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"dl_out_mask\" -q sc2mac_dat_b_mask");
//: my $i;
//: for($i = 0; $i < 64; $i ++) {
//: &eperl::flop("-wid 8 -norst -en \"dl_out_mask[${i}]\" -d \"dl_out_data${i}\" -q sc2mac_dat_a_data${i}");
//: }
//: print "\n\n";
//:
//: for($i = 0; $i < 64; $i ++) {
//: &eperl::flop("-wid 8  -norst -en \"dl_out_mask[${i}]\" -d \"dl_out_data${i}\" -q sc2mac_dat_b_data${i}");
//: }
//: print "\n\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_pvld_d1 <= 1'b0;
   end else begin
       dl_out_pvld_d1 <= dl_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_a_pvld <= 1'b0;
   end else begin
       sc2mac_dat_a_pvld <= dl_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_b_pvld <= 1'b0;
   end else begin
       sc2mac_dat_b_pvld <= dl_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_a_pd <= {9{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_a_pd <= sc2mac_dat_pd_w;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_a_pd <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_b_pd <= {9{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_b_pd <= sc2mac_dat_pd_w;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_b_pd <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_a_mask <= {64{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_a_mask <= dl_out_mask;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_a_mask <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_b_mask <= {64{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_b_mask <= dl_out_mask;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_b_mask <= 'bx;
       // VCS coverage on
       end
   end
end
reg [7:0] sc2mac_dat_a_data0;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[0]) == 1'b1) begin
           sc2mac_dat_a_data0 <= dl_out_data0;
       // VCS coverage off
       end else if ((dl_out_mask[0]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data0 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data1;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[1]) == 1'b1) begin
           sc2mac_dat_a_data1 <= dl_out_data1;
       // VCS coverage off
       end else if ((dl_out_mask[1]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data1 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data2;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[2]) == 1'b1) begin
           sc2mac_dat_a_data2 <= dl_out_data2;
       // VCS coverage off
       end else if ((dl_out_mask[2]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data2 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data3;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[3]) == 1'b1) begin
           sc2mac_dat_a_data3 <= dl_out_data3;
       // VCS coverage off
       end else if ((dl_out_mask[3]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data3 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data4;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[4]) == 1'b1) begin
           sc2mac_dat_a_data4 <= dl_out_data4;
       // VCS coverage off
       end else if ((dl_out_mask[4]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data4 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data5;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[5]) == 1'b1) begin
           sc2mac_dat_a_data5 <= dl_out_data5;
       // VCS coverage off
       end else if ((dl_out_mask[5]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data5 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data6;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[6]) == 1'b1) begin
           sc2mac_dat_a_data6 <= dl_out_data6;
       // VCS coverage off
       end else if ((dl_out_mask[6]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data6 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data7;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[7]) == 1'b1) begin
           sc2mac_dat_a_data7 <= dl_out_data7;
       // VCS coverage off
       end else if ((dl_out_mask[7]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data7 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data8;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[8]) == 1'b1) begin
           sc2mac_dat_a_data8 <= dl_out_data8;
       // VCS coverage off
       end else if ((dl_out_mask[8]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data8 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data9;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[9]) == 1'b1) begin
           sc2mac_dat_a_data9 <= dl_out_data9;
       // VCS coverage off
       end else if ((dl_out_mask[9]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data9 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data10;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[10]) == 1'b1) begin
           sc2mac_dat_a_data10 <= dl_out_data10;
       // VCS coverage off
       end else if ((dl_out_mask[10]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data10 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data11;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[11]) == 1'b1) begin
           sc2mac_dat_a_data11 <= dl_out_data11;
       // VCS coverage off
       end else if ((dl_out_mask[11]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data11 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data12;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[12]) == 1'b1) begin
           sc2mac_dat_a_data12 <= dl_out_data12;
       // VCS coverage off
       end else if ((dl_out_mask[12]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data12 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data13;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[13]) == 1'b1) begin
           sc2mac_dat_a_data13 <= dl_out_data13;
       // VCS coverage off
       end else if ((dl_out_mask[13]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data13 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data14;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[14]) == 1'b1) begin
           sc2mac_dat_a_data14 <= dl_out_data14;
       // VCS coverage off
       end else if ((dl_out_mask[14]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data14 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data15;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[15]) == 1'b1) begin
           sc2mac_dat_a_data15 <= dl_out_data15;
       // VCS coverage off
       end else if ((dl_out_mask[15]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data15 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data16;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[16]) == 1'b1) begin
           sc2mac_dat_a_data16 <= dl_out_data16;
       // VCS coverage off
       end else if ((dl_out_mask[16]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data16 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data17;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[17]) == 1'b1) begin
           sc2mac_dat_a_data17 <= dl_out_data17;
       // VCS coverage off
       end else if ((dl_out_mask[17]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data17 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data18;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[18]) == 1'b1) begin
           sc2mac_dat_a_data18 <= dl_out_data18;
       // VCS coverage off
       end else if ((dl_out_mask[18]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data18 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data19;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[19]) == 1'b1) begin
           sc2mac_dat_a_data19 <= dl_out_data19;
       // VCS coverage off
       end else if ((dl_out_mask[19]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data19 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data20;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[20]) == 1'b1) begin
           sc2mac_dat_a_data20 <= dl_out_data20;
       // VCS coverage off
       end else if ((dl_out_mask[20]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data20 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data21;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[21]) == 1'b1) begin
           sc2mac_dat_a_data21 <= dl_out_data21;
       // VCS coverage off
       end else if ((dl_out_mask[21]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data21 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data22;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[22]) == 1'b1) begin
           sc2mac_dat_a_data22 <= dl_out_data22;
       // VCS coverage off
       end else if ((dl_out_mask[22]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data22 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data23;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[23]) == 1'b1) begin
           sc2mac_dat_a_data23 <= dl_out_data23;
       // VCS coverage off
       end else if ((dl_out_mask[23]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data23 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data24;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[24]) == 1'b1) begin
           sc2mac_dat_a_data24 <= dl_out_data24;
       // VCS coverage off
       end else if ((dl_out_mask[24]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data24 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data25;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[25]) == 1'b1) begin
           sc2mac_dat_a_data25 <= dl_out_data25;
       // VCS coverage off
       end else if ((dl_out_mask[25]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data25 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data26;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[26]) == 1'b1) begin
           sc2mac_dat_a_data26 <= dl_out_data26;
       // VCS coverage off
       end else if ((dl_out_mask[26]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data26 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data27;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[27]) == 1'b1) begin
           sc2mac_dat_a_data27 <= dl_out_data27;
       // VCS coverage off
       end else if ((dl_out_mask[27]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data27 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data28;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[28]) == 1'b1) begin
           sc2mac_dat_a_data28 <= dl_out_data28;
       // VCS coverage off
       end else if ((dl_out_mask[28]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data28 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data29;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[29]) == 1'b1) begin
           sc2mac_dat_a_data29 <= dl_out_data29;
       // VCS coverage off
       end else if ((dl_out_mask[29]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data29 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data30;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[30]) == 1'b1) begin
           sc2mac_dat_a_data30 <= dl_out_data30;
       // VCS coverage off
       end else if ((dl_out_mask[30]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data30 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data31;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[31]) == 1'b1) begin
           sc2mac_dat_a_data31 <= dl_out_data31;
       // VCS coverage off
       end else if ((dl_out_mask[31]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data31 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data32;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[32]) == 1'b1) begin
           sc2mac_dat_a_data32 <= dl_out_data32;
       // VCS coverage off
       end else if ((dl_out_mask[32]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data32 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data33;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[33]) == 1'b1) begin
           sc2mac_dat_a_data33 <= dl_out_data33;
       // VCS coverage off
       end else if ((dl_out_mask[33]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data33 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data34;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[34]) == 1'b1) begin
           sc2mac_dat_a_data34 <= dl_out_data34;
       // VCS coverage off
       end else if ((dl_out_mask[34]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data34 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data35;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[35]) == 1'b1) begin
           sc2mac_dat_a_data35 <= dl_out_data35;
       // VCS coverage off
       end else if ((dl_out_mask[35]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data35 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data36;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[36]) == 1'b1) begin
           sc2mac_dat_a_data36 <= dl_out_data36;
       // VCS coverage off
       end else if ((dl_out_mask[36]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data36 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data37;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[37]) == 1'b1) begin
           sc2mac_dat_a_data37 <= dl_out_data37;
       // VCS coverage off
       end else if ((dl_out_mask[37]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data37 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data38;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[38]) == 1'b1) begin
           sc2mac_dat_a_data38 <= dl_out_data38;
       // VCS coverage off
       end else if ((dl_out_mask[38]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data38 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data39;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[39]) == 1'b1) begin
           sc2mac_dat_a_data39 <= dl_out_data39;
       // VCS coverage off
       end else if ((dl_out_mask[39]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data39 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data40;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[40]) == 1'b1) begin
           sc2mac_dat_a_data40 <= dl_out_data40;
       // VCS coverage off
       end else if ((dl_out_mask[40]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data40 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data41;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[41]) == 1'b1) begin
           sc2mac_dat_a_data41 <= dl_out_data41;
       // VCS coverage off
       end else if ((dl_out_mask[41]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data41 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data42;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[42]) == 1'b1) begin
           sc2mac_dat_a_data42 <= dl_out_data42;
       // VCS coverage off
       end else if ((dl_out_mask[42]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data42 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data43;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[43]) == 1'b1) begin
           sc2mac_dat_a_data43 <= dl_out_data43;
       // VCS coverage off
       end else if ((dl_out_mask[43]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data43 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data44;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[44]) == 1'b1) begin
           sc2mac_dat_a_data44 <= dl_out_data44;
       // VCS coverage off
       end else if ((dl_out_mask[44]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data44 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data45;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[45]) == 1'b1) begin
           sc2mac_dat_a_data45 <= dl_out_data45;
       // VCS coverage off
       end else if ((dl_out_mask[45]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data45 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data46;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[46]) == 1'b1) begin
           sc2mac_dat_a_data46 <= dl_out_data46;
       // VCS coverage off
       end else if ((dl_out_mask[46]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data46 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data47;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[47]) == 1'b1) begin
           sc2mac_dat_a_data47 <= dl_out_data47;
       // VCS coverage off
       end else if ((dl_out_mask[47]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data47 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data48;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[48]) == 1'b1) begin
           sc2mac_dat_a_data48 <= dl_out_data48;
       // VCS coverage off
       end else if ((dl_out_mask[48]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data48 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data49;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[49]) == 1'b1) begin
           sc2mac_dat_a_data49 <= dl_out_data49;
       // VCS coverage off
       end else if ((dl_out_mask[49]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data49 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data50;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[50]) == 1'b1) begin
           sc2mac_dat_a_data50 <= dl_out_data50;
       // VCS coverage off
       end else if ((dl_out_mask[50]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data50 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data51;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[51]) == 1'b1) begin
           sc2mac_dat_a_data51 <= dl_out_data51;
       // VCS coverage off
       end else if ((dl_out_mask[51]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data51 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data52;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[52]) == 1'b1) begin
           sc2mac_dat_a_data52 <= dl_out_data52;
       // VCS coverage off
       end else if ((dl_out_mask[52]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data52 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data53;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[53]) == 1'b1) begin
           sc2mac_dat_a_data53 <= dl_out_data53;
       // VCS coverage off
       end else if ((dl_out_mask[53]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data53 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data54;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[54]) == 1'b1) begin
           sc2mac_dat_a_data54 <= dl_out_data54;
       // VCS coverage off
       end else if ((dl_out_mask[54]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data54 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data55;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[55]) == 1'b1) begin
           sc2mac_dat_a_data55 <= dl_out_data55;
       // VCS coverage off
       end else if ((dl_out_mask[55]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data55 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data56;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[56]) == 1'b1) begin
           sc2mac_dat_a_data56 <= dl_out_data56;
       // VCS coverage off
       end else if ((dl_out_mask[56]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data56 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data57;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[57]) == 1'b1) begin
           sc2mac_dat_a_data57 <= dl_out_data57;
       // VCS coverage off
       end else if ((dl_out_mask[57]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data57 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data58;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[58]) == 1'b1) begin
           sc2mac_dat_a_data58 <= dl_out_data58;
       // VCS coverage off
       end else if ((dl_out_mask[58]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data58 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data59;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[59]) == 1'b1) begin
           sc2mac_dat_a_data59 <= dl_out_data59;
       // VCS coverage off
       end else if ((dl_out_mask[59]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data59 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data60;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[60]) == 1'b1) begin
           sc2mac_dat_a_data60 <= dl_out_data60;
       // VCS coverage off
       end else if ((dl_out_mask[60]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data60 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data61;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[61]) == 1'b1) begin
           sc2mac_dat_a_data61 <= dl_out_data61;
       // VCS coverage off
       end else if ((dl_out_mask[61]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data61 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data62;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[62]) == 1'b1) begin
           sc2mac_dat_a_data62 <= dl_out_data62;
       // VCS coverage off
       end else if ((dl_out_mask[62]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data62 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data63;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[63]) == 1'b1) begin
           sc2mac_dat_a_data63 <= dl_out_data63;
       // VCS coverage off
       end else if ((dl_out_mask[63]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data63 <= 'bx;
       // VCS coverage on
       end
end


reg [7:0] sc2mac_dat_b_data0;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[0]) == 1'b1) begin
           sc2mac_dat_b_data0 <= dl_out_data0;
       // VCS coverage off
       end else if ((dl_out_mask[0]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data0 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data1;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[1]) == 1'b1) begin
           sc2mac_dat_b_data1 <= dl_out_data1;
       // VCS coverage off
       end else if ((dl_out_mask[1]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data1 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data2;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[2]) == 1'b1) begin
           sc2mac_dat_b_data2 <= dl_out_data2;
       // VCS coverage off
       end else if ((dl_out_mask[2]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data2 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data3;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[3]) == 1'b1) begin
           sc2mac_dat_b_data3 <= dl_out_data3;
       // VCS coverage off
       end else if ((dl_out_mask[3]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data3 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data4;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[4]) == 1'b1) begin
           sc2mac_dat_b_data4 <= dl_out_data4;
       // VCS coverage off
       end else if ((dl_out_mask[4]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data4 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data5;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[5]) == 1'b1) begin
           sc2mac_dat_b_data5 <= dl_out_data5;
       // VCS coverage off
       end else if ((dl_out_mask[5]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data5 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data6;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[6]) == 1'b1) begin
           sc2mac_dat_b_data6 <= dl_out_data6;
       // VCS coverage off
       end else if ((dl_out_mask[6]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data6 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data7;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[7]) == 1'b1) begin
           sc2mac_dat_b_data7 <= dl_out_data7;
       // VCS coverage off
       end else if ((dl_out_mask[7]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data7 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data8;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[8]) == 1'b1) begin
           sc2mac_dat_b_data8 <= dl_out_data8;
       // VCS coverage off
       end else if ((dl_out_mask[8]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data8 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data9;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[9]) == 1'b1) begin
           sc2mac_dat_b_data9 <= dl_out_data9;
       // VCS coverage off
       end else if ((dl_out_mask[9]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data9 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data10;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[10]) == 1'b1) begin
           sc2mac_dat_b_data10 <= dl_out_data10;
       // VCS coverage off
       end else if ((dl_out_mask[10]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data10 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data11;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[11]) == 1'b1) begin
           sc2mac_dat_b_data11 <= dl_out_data11;
       // VCS coverage off
       end else if ((dl_out_mask[11]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data11 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data12;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[12]) == 1'b1) begin
           sc2mac_dat_b_data12 <= dl_out_data12;
       // VCS coverage off
       end else if ((dl_out_mask[12]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data12 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data13;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[13]) == 1'b1) begin
           sc2mac_dat_b_data13 <= dl_out_data13;
       // VCS coverage off
       end else if ((dl_out_mask[13]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data13 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data14;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[14]) == 1'b1) begin
           sc2mac_dat_b_data14 <= dl_out_data14;
       // VCS coverage off
       end else if ((dl_out_mask[14]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data14 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data15;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[15]) == 1'b1) begin
           sc2mac_dat_b_data15 <= dl_out_data15;
       // VCS coverage off
       end else if ((dl_out_mask[15]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data15 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data16;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[16]) == 1'b1) begin
           sc2mac_dat_b_data16 <= dl_out_data16;
       // VCS coverage off
       end else if ((dl_out_mask[16]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data16 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data17;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[17]) == 1'b1) begin
           sc2mac_dat_b_data17 <= dl_out_data17;
       // VCS coverage off
       end else if ((dl_out_mask[17]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data17 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data18;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[18]) == 1'b1) begin
           sc2mac_dat_b_data18 <= dl_out_data18;
       // VCS coverage off
       end else if ((dl_out_mask[18]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data18 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data19;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[19]) == 1'b1) begin
           sc2mac_dat_b_data19 <= dl_out_data19;
       // VCS coverage off
       end else if ((dl_out_mask[19]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data19 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data20;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[20]) == 1'b1) begin
           sc2mac_dat_b_data20 <= dl_out_data20;
       // VCS coverage off
       end else if ((dl_out_mask[20]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data20 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data21;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[21]) == 1'b1) begin
           sc2mac_dat_b_data21 <= dl_out_data21;
       // VCS coverage off
       end else if ((dl_out_mask[21]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data21 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data22;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[22]) == 1'b1) begin
           sc2mac_dat_b_data22 <= dl_out_data22;
       // VCS coverage off
       end else if ((dl_out_mask[22]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data22 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data23;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[23]) == 1'b1) begin
           sc2mac_dat_b_data23 <= dl_out_data23;
       // VCS coverage off
       end else if ((dl_out_mask[23]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data23 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data24;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[24]) == 1'b1) begin
           sc2mac_dat_b_data24 <= dl_out_data24;
       // VCS coverage off
       end else if ((dl_out_mask[24]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data24 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data25;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[25]) == 1'b1) begin
           sc2mac_dat_b_data25 <= dl_out_data25;
       // VCS coverage off
       end else if ((dl_out_mask[25]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data25 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data26;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[26]) == 1'b1) begin
           sc2mac_dat_b_data26 <= dl_out_data26;
       // VCS coverage off
       end else if ((dl_out_mask[26]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data26 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data27;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[27]) == 1'b1) begin
           sc2mac_dat_b_data27 <= dl_out_data27;
       // VCS coverage off
       end else if ((dl_out_mask[27]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data27 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data28;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[28]) == 1'b1) begin
           sc2mac_dat_b_data28 <= dl_out_data28;
       // VCS coverage off
       end else if ((dl_out_mask[28]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data28 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data29;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[29]) == 1'b1) begin
           sc2mac_dat_b_data29 <= dl_out_data29;
       // VCS coverage off
       end else if ((dl_out_mask[29]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data29 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data30;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[30]) == 1'b1) begin
           sc2mac_dat_b_data30 <= dl_out_data30;
       // VCS coverage off
       end else if ((dl_out_mask[30]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data30 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data31;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[31]) == 1'b1) begin
           sc2mac_dat_b_data31 <= dl_out_data31;
       // VCS coverage off
       end else if ((dl_out_mask[31]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data31 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data32;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[32]) == 1'b1) begin
           sc2mac_dat_b_data32 <= dl_out_data32;
       // VCS coverage off
       end else if ((dl_out_mask[32]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data32 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data33;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[33]) == 1'b1) begin
           sc2mac_dat_b_data33 <= dl_out_data33;
       // VCS coverage off
       end else if ((dl_out_mask[33]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data33 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data34;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[34]) == 1'b1) begin
           sc2mac_dat_b_data34 <= dl_out_data34;
       // VCS coverage off
       end else if ((dl_out_mask[34]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data34 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data35;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[35]) == 1'b1) begin
           sc2mac_dat_b_data35 <= dl_out_data35;
       // VCS coverage off
       end else if ((dl_out_mask[35]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data35 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data36;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[36]) == 1'b1) begin
           sc2mac_dat_b_data36 <= dl_out_data36;
       // VCS coverage off
       end else if ((dl_out_mask[36]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data36 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data37;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[37]) == 1'b1) begin
           sc2mac_dat_b_data37 <= dl_out_data37;
       // VCS coverage off
       end else if ((dl_out_mask[37]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data37 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data38;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[38]) == 1'b1) begin
           sc2mac_dat_b_data38 <= dl_out_data38;
       // VCS coverage off
       end else if ((dl_out_mask[38]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data38 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data39;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[39]) == 1'b1) begin
           sc2mac_dat_b_data39 <= dl_out_data39;
       // VCS coverage off
       end else if ((dl_out_mask[39]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data39 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data40;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[40]) == 1'b1) begin
           sc2mac_dat_b_data40 <= dl_out_data40;
       // VCS coverage off
       end else if ((dl_out_mask[40]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data40 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data41;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[41]) == 1'b1) begin
           sc2mac_dat_b_data41 <= dl_out_data41;
       // VCS coverage off
       end else if ((dl_out_mask[41]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data41 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data42;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[42]) == 1'b1) begin
           sc2mac_dat_b_data42 <= dl_out_data42;
       // VCS coverage off
       end else if ((dl_out_mask[42]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data42 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data43;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[43]) == 1'b1) begin
           sc2mac_dat_b_data43 <= dl_out_data43;
       // VCS coverage off
       end else if ((dl_out_mask[43]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data43 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data44;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[44]) == 1'b1) begin
           sc2mac_dat_b_data44 <= dl_out_data44;
       // VCS coverage off
       end else if ((dl_out_mask[44]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data44 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data45;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[45]) == 1'b1) begin
           sc2mac_dat_b_data45 <= dl_out_data45;
       // VCS coverage off
       end else if ((dl_out_mask[45]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data45 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data46;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[46]) == 1'b1) begin
           sc2mac_dat_b_data46 <= dl_out_data46;
       // VCS coverage off
       end else if ((dl_out_mask[46]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data46 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data47;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[47]) == 1'b1) begin
           sc2mac_dat_b_data47 <= dl_out_data47;
       // VCS coverage off
       end else if ((dl_out_mask[47]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data47 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data48;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[48]) == 1'b1) begin
           sc2mac_dat_b_data48 <= dl_out_data48;
       // VCS coverage off
       end else if ((dl_out_mask[48]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data48 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data49;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[49]) == 1'b1) begin
           sc2mac_dat_b_data49 <= dl_out_data49;
       // VCS coverage off
       end else if ((dl_out_mask[49]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data49 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data50;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[50]) == 1'b1) begin
           sc2mac_dat_b_data50 <= dl_out_data50;
       // VCS coverage off
       end else if ((dl_out_mask[50]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data50 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data51;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[51]) == 1'b1) begin
           sc2mac_dat_b_data51 <= dl_out_data51;
       // VCS coverage off
       end else if ((dl_out_mask[51]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data51 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data52;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[52]) == 1'b1) begin
           sc2mac_dat_b_data52 <= dl_out_data52;
       // VCS coverage off
       end else if ((dl_out_mask[52]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data52 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data53;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[53]) == 1'b1) begin
           sc2mac_dat_b_data53 <= dl_out_data53;
       // VCS coverage off
       end else if ((dl_out_mask[53]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data53 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data54;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[54]) == 1'b1) begin
           sc2mac_dat_b_data54 <= dl_out_data54;
       // VCS coverage off
       end else if ((dl_out_mask[54]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data54 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data55;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[55]) == 1'b1) begin
           sc2mac_dat_b_data55 <= dl_out_data55;
       // VCS coverage off
       end else if ((dl_out_mask[55]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data55 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data56;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[56]) == 1'b1) begin
           sc2mac_dat_b_data56 <= dl_out_data56;
       // VCS coverage off
       end else if ((dl_out_mask[56]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data56 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data57;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[57]) == 1'b1) begin
           sc2mac_dat_b_data57 <= dl_out_data57;
       // VCS coverage off
       end else if ((dl_out_mask[57]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data57 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data58;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[58]) == 1'b1) begin
           sc2mac_dat_b_data58 <= dl_out_data58;
       // VCS coverage off
       end else if ((dl_out_mask[58]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data58 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data59;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[59]) == 1'b1) begin
           sc2mac_dat_b_data59 <= dl_out_data59;
       // VCS coverage off
       end else if ((dl_out_mask[59]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data59 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data60;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[60]) == 1'b1) begin
           sc2mac_dat_b_data60 <= dl_out_data60;
       // VCS coverage off
       end else if ((dl_out_mask[60]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data60 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data61;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[61]) == 1'b1) begin
           sc2mac_dat_b_data61 <= dl_out_data61;
       // VCS coverage off
       end else if ((dl_out_mask[61]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data61 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data62;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[62]) == 1'b1) begin
           sc2mac_dat_b_data62 <= dl_out_data62;
       // VCS coverage off
       end else if ((dl_out_mask[62]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data62 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data63;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[63]) == 1'b1) begin
           sc2mac_dat_b_data63 <= dl_out_data63;
       // VCS coverage off
       end else if ((dl_out_mask[63]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data63 <= 'bx;
       // VCS coverage on
       end
end


endmodule // NV_NVDLA_CSC_dl

module NV_soDLA_CSC_dl_for_check( // @[:@3.2]
  input          io_nvdla_core_clk, // @[:@6.4]
  input          io_nvdla_core_ng_clk, // @[:@6.4]
  input          io_nvdla_core_rstn, // @[:@6.4]
  input  [1:0]   io_sc_state, // @[:@6.4]
  input          io_sg2dl_pd_valid, // @[:@6.4]
  input  [30:0]  io_sg2dl_pd_bits, // @[:@6.4]
  input          io_sg2dl_reuse_rls, // @[:@6.4]
  input          io_cdma2sc_dat_updt_valid, // @[:@6.4]
  input  [14:0]  io_cdma2sc_dat_updt_bits_entries, // @[:@6.4]
  input  [13:0]  io_cdma2sc_dat_updt_bits_slices, // @[:@6.4]
  input          io_sc2cdma_dat_pending_req, // @[:@6.4]
  output         io_sc2cdma_dat_updt_valid, // @[:@6.4]
  output [14:0]  io_sc2cdma_dat_updt_bits_entries, // @[:@6.4]
  output [13:0]  io_sc2cdma_dat_updt_bits_slices, // @[:@6.4]
  output         io_sc2buf_dat_rd_addr_valid, // @[:@6.4]
  output [12:0]  io_sc2buf_dat_rd_addr_bits, // @[:@6.4]
  input          io_sc2buf_dat_rd_data_valid, // @[:@6.4]
  input  [511:0] io_sc2buf_dat_rd_data_bits, // @[:@6.4]
  output         io_sc2mac_dat_a_valid, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_0, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_1, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_2, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_3, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_4, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_5, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_6, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_7, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_8, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_9, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_10, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_11, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_12, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_13, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_14, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_15, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_16, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_17, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_18, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_19, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_20, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_21, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_22, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_23, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_24, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_25, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_26, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_27, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_28, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_29, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_30, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_31, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_32, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_33, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_34, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_35, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_36, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_37, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_38, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_39, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_40, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_41, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_42, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_43, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_44, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_45, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_46, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_47, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_48, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_49, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_50, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_51, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_52, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_53, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_54, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_55, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_56, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_57, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_58, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_59, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_60, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_61, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_62, // @[:@6.4]
  output         io_sc2mac_dat_a_bits_mask_63, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_0, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_1, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_2, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_3, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_4, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_5, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_6, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_7, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_8, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_9, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_10, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_11, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_12, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_13, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_14, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_15, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_16, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_17, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_18, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_19, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_20, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_21, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_22, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_23, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_24, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_25, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_26, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_27, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_28, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_29, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_30, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_31, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_32, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_33, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_34, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_35, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_36, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_37, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_38, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_39, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_40, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_41, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_42, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_43, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_44, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_45, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_46, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_47, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_48, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_49, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_50, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_51, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_52, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_53, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_54, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_55, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_56, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_57, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_58, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_59, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_60, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_61, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_62, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_bits_data_63, // @[:@6.4]
  output [8:0]   io_sc2mac_dat_a_bits_pd, // @[:@6.4]
  output         io_sc2mac_dat_b_valid, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_0, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_1, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_2, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_3, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_4, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_5, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_6, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_7, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_8, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_9, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_10, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_11, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_12, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_13, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_14, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_15, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_16, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_17, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_18, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_19, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_20, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_21, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_22, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_23, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_24, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_25, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_26, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_27, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_28, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_29, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_30, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_31, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_32, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_33, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_34, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_35, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_36, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_37, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_38, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_39, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_40, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_41, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_42, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_43, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_44, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_45, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_46, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_47, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_48, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_49, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_50, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_51, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_52, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_53, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_54, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_55, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_56, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_57, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_58, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_59, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_60, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_61, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_62, // @[:@6.4]
  output         io_sc2mac_dat_b_bits_mask_63, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_0, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_1, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_2, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_3, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_4, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_5, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_6, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_7, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_8, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_9, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_10, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_11, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_12, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_13, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_14, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_15, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_16, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_17, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_18, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_19, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_20, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_21, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_22, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_23, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_24, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_25, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_26, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_27, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_28, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_29, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_30, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_31, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_32, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_33, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_34, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_35, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_36, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_37, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_38, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_39, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_40, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_41, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_42, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_43, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_44, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_45, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_46, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_47, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_48, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_49, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_50, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_51, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_52, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_53, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_54, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_55, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_56, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_57, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_58, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_59, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_60, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_61, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_62, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_bits_data_63, // @[:@6.4]
  output [8:0]   io_sc2mac_dat_b_bits_pd, // @[:@6.4]
  input          io_reg2dp_op_en, // @[:@6.4]
  input          io_reg2dp_conv_mode, // @[:@6.4]
  input  [4:0]   io_reg2dp_batches, // @[:@6.4]
  input  [1:0]   io_reg2dp_proc_precision, // @[:@6.4]
  input          io_reg2dp_datain_format, // @[:@6.4]
  input          io_reg2dp_skip_data_rls, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_channel_ext, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_height_ext, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_width_ext, // @[:@6.4]
  input  [1:0]   io_reg2dp_y_extension, // @[:@6.4]
  input  [12:0]  io_reg2dp_weight_channel_ext, // @[:@6.4]
  input  [13:0]  io_reg2dp_entries, // @[:@6.4]
  input  [12:0]  io_reg2dp_dataout_width, // @[:@6.4]
  input  [11:0]  io_reg2dp_rls_slices, // @[:@6.4]
  input  [2:0]   io_reg2dp_conv_x_stride_ext, // @[:@6.4]
  input  [2:0]   io_reg2dp_conv_y_stride_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_x_dilation_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_y_dilation_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_pad_left, // @[:@6.4]
  input  [4:0]   io_reg2dp_pad_top, // @[:@6.4]
  input  [15:0]  io_reg2dp_pad_value, // @[:@6.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@6.4]
  input  [1:0]   io_reg2dp_pra_truncate, // @[:@6.4]
  output         io_slcg_wg_en // @[:@6.4]
);
  wire  _T_623; // @[NV_NVDLA_CSC_dl_for_check.scala 73:38:@8.4]
  wire  _T_625; // @[NV_NVDLA_CSC_dl_for_check.scala 77:31:@9.4]
  wire  _T_629; // @[NV_NVDLA_CSC_dl_for_check.scala 79:31:@11.4]
  wire  _T_633; // @[NV_NVDLA_CSC_dl_for_check.scala 86:32:@14.4]
  wire  _T_637; // @[NV_NVDLA_CSC_dl_for_check.scala 88:35:@16.4]
  wire  _T_638; // @[NV_NVDLA_CSC_dl_for_check.scala 89:22:@17.4]
  wire [6:0] _T_643; // @[NV_NVDLA_CSC_dl_for_check.scala 96:53:@18.4]
  wire [6:0] _T_645; // @[NV_NVDLA_CSC_dl_for_check.scala 96:24:@19.4]
  wire [2:0] _T_646; // @[NV_NVDLA_CSC_dl_for_check.scala 96:100:@20.4]
  wire [2:0] _T_648; // @[NV_NVDLA_CSC_dl_for_check.scala 97:22:@21.4]
  wire [3:0] _T_650; // @[NV_NVDLA_CSC_dl_for_check.scala 98:34:@22.4]
  wire [3:0] _T_651; // @[NV_NVDLA_CSC_dl_for_check.scala 98:34:@23.4]
  wire [3:0] _T_653; // @[NV_NVDLA_CSC_dl_for_check.scala 99:51:@24.4]
  wire [1:0] _T_654; // @[NV_NVDLA_CSC_dl_for_check.scala 100:62:@25.4]
  wire [5:0] _T_657; // @[Cat.scala 30:58:@26.4]
  wire [4:0] _T_660; // @[Cat.scala 30:58:@27.4]
  wire [4:0] _GEN_671; // @[NV_NVDLA_CSC_dl_for_check.scala 102:74:@28.4]
  wire [5:0] _T_661; // @[NV_NVDLA_CSC_dl_for_check.scala 102:74:@28.4]
  wire  _T_662; // @[Mux.scala 46:19:@29.4]
  wire [5:0] _T_663; // @[Mux.scala 46:16:@30.4]
  wire  _T_664; // @[Mux.scala 46:19:@31.4]
  wire [5:0] _T_665; // @[Mux.scala 46:16:@32.4]
  wire  _T_667; // @[NV_NVDLA_CSC_dl_for_check.scala 104:88:@33.4]
  wire [5:0] _T_673; // @[NV_NVDLA_CSC_dl_for_check.scala 104:172:@35.4]
  wire [5:0] _T_674; // @[NV_NVDLA_CSC_dl_for_check.scala 104:58:@36.4]
  wire [6:0] _T_677; // @[Cat.scala 30:58:@37.4]
  wire [6:0] _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 105:81:@38.4]
  wire [7:0] _T_678; // @[NV_NVDLA_CSC_dl_for_check.scala 105:81:@38.4]
  wire [6:0] _T_679; // @[NV_NVDLA_CSC_dl_for_check.scala 105:81:@39.4]
  wire [6:0] _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@41.4]
  wire [7:0] _T_681; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@41.4]
  wire [6:0] _T_682; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@42.4]
  wire [6:0] _T_685; // @[NV_NVDLA_CSC_dl_for_check.scala 106:58:@44.4]
  wire [5:0] _T_686; // @[NV_NVDLA_CSC_dl_for_check.scala 106:58:@45.4]
  wire  _T_687; // @[Mux.scala 46:19:@46.4]
  wire [5:0] _T_688; // @[Mux.scala 46:16:@47.4]
  wire  _T_689; // @[Mux.scala 46:19:@48.4]
  wire [6:0] _T_690; // @[Mux.scala 46:16:@49.4]
  wire [6:0] _T_693; // @[NV_NVDLA_CSC_dl_for_check.scala 107:80:@51.4]
  wire [7:0] _T_696; // @[Cat.scala 30:58:@52.4]
  wire [6:0] _T_701; // @[Mux.scala 46:16:@55.4]
  wire [7:0] _T_703; // @[Mux.scala 46:16:@57.4]
  wire [11:0] _T_705; // @[Cat.scala 30:58:@58.4]
  wire [3:0] _T_707; // @[NV_NVDLA_CSC_dl_for_check.scala 117:52:@59.4]
  wire [5:0] _T_710; // @[NV_NVDLA_CSC_dl_for_check.scala 118:60:@60.4]
  wire [5:0] _T_711; // @[NV_NVDLA_CSC_dl_for_check.scala 118:21:@61.4]
  wire [5:0] _T_714; // @[NV_NVDLA_CSC_dl_for_check.scala 119:60:@62.4]
  wire [5:0] _T_715; // @[NV_NVDLA_CSC_dl_for_check.scala 119:21:@63.4]
  reg  _T_718; // @[NV_NVDLA_CSC_dl_for_check.scala 121:26:@64.4]
  reg [31:0] _RAND_0;
  reg [5:0] _T_725; // @[NV_NVDLA_CSC_dl_for_check.scala 122:25:@66.4]
  reg [31:0] _RAND_1;
  reg [13:0] _T_732; // @[NV_NVDLA_CSC_dl_for_check.scala 123:25:@68.4]
  reg [31:0] _RAND_2;
  reg [13:0] _T_739; // @[NV_NVDLA_CSC_dl_for_check.scala 124:29:@70.4]
  reg [31:0] _RAND_3;
  reg [14:0] _T_746; // @[NV_NVDLA_CSC_dl_for_check.scala 125:22:@72.4]
  reg [31:0] _RAND_4;
  reg [14:0] _T_753; // @[NV_NVDLA_CSC_dl_for_check.scala 126:28:@74.4]
  reg [31:0] _RAND_5;
  reg [12:0] _T_760; // @[NV_NVDLA_CSC_dl_for_check.scala 127:32:@76.4]
  reg [31:0] _RAND_6;
  reg [14:0] _T_774; // @[NV_NVDLA_CSC_dl_for_check.scala 129:26:@80.4]
  reg [31:0] _RAND_7;
  reg [11:0] _T_781; // @[NV_NVDLA_CSC_dl_for_check.scala 130:30:@82.4]
  reg [31:0] _RAND_8;
  reg [11:0] _T_788; // @[NV_NVDLA_CSC_dl_for_check.scala 131:30:@84.4]
  reg [31:0] _RAND_9;
  reg [13:0] _T_795; // @[NV_NVDLA_CSC_dl_for_check.scala 132:25:@86.4]
  reg [31:0] _RAND_10;
  wire [14:0] _T_797; // @[NV_NVDLA_CSC_dl_for_check.scala 135:43:@87.4]
  wire [20:0] _T_799; // @[NV_NVDLA_CSC_dl_for_check.scala 136:41:@89.4]
  wire [14:0] _T_800; // @[NV_NVDLA_CSC_dl_for_check.scala 136:56:@90.4]
  wire [11:0] _T_801; // @[NV_NVDLA_CSC_dl_for_check.scala 138:37:@91.4]
  wire [14:0] _GEN_674; // @[NV_NVDLA_CSC_dl_for_check.scala 139:34:@92.4]
  wire [20:0] _T_802; // @[NV_NVDLA_CSC_dl_for_check.scala 139:34:@92.4]
  wire [11:0] _T_803; // @[NV_NVDLA_CSC_dl_for_check.scala 139:47:@93.4]
  wire [14:0] _GEN_675; // @[NV_NVDLA_CSC_dl_for_check.scala 140:34:@94.4]
  wire [28:0] _T_804; // @[NV_NVDLA_CSC_dl_for_check.scala 140:34:@94.4]
  wire [11:0] _T_805; // @[NV_NVDLA_CSC_dl_for_check.scala 140:51:@95.4]
  wire [12:0] _T_807; // @[NV_NVDLA_CSC_dl_for_check.scala 141:41:@96.4]
  wire [11:0] _T_808; // @[NV_NVDLA_CSC_dl_for_check.scala 141:41:@97.4]
  wire [13:0] _T_810; // @[NV_NVDLA_CSC_dl_for_check.scala 142:77:@98.4]
  wire [12:0] _GEN_676; // @[NV_NVDLA_CSC_dl_for_check.scala 142:113:@99.4]
  wire [13:0] _T_811; // @[NV_NVDLA_CSC_dl_for_check.scala 142:113:@99.4]
  wire [13:0] _T_812; // @[NV_NVDLA_CSC_dl_for_check.scala 142:113:@100.4]
  wire [13:0] _T_813; // @[NV_NVDLA_CSC_dl_for_check.scala 142:23:@101.4]
  wire [13:0] _T_814; // @[NV_NVDLA_CSC_dl_for_check.scala 143:24:@102.4]
  wire [14:0] _GEN_677; // @[NV_NVDLA_CSC_dl_for_check.scala 144:38:@103.4]
  wire [28:0] _T_815; // @[NV_NVDLA_CSC_dl_for_check.scala 144:38:@103.4]
  wire [14:0] _T_816; // @[NV_NVDLA_CSC_dl_for_check.scala 144:54:@104.4]
  reg [33:0] _T_834; // @[NV_NVDLA_CSC_dl_for_check.scala 149:24:@110.4]
  reg [63:0] _RAND_11;
  reg [4:0] _T_841; // @[NV_NVDLA_CSC_dl_for_check.scala 150:24:@112.4]
  reg [31:0] _RAND_12;
  reg [13:0] _T_848; // @[NV_NVDLA_CSC_dl_for_check.scala 151:27:@114.4]
  reg [31:0] _RAND_13;
  reg [12:0] _T_855; // @[NV_NVDLA_CSC_dl_for_check.scala 152:31:@116.4]
  reg [31:0] _RAND_14;
  reg [12:0] _T_862; // @[NV_NVDLA_CSC_dl_for_check.scala 153:32:@118.4]
  reg [31:0] _RAND_15;
  reg [10:0] _T_869; // @[NV_NVDLA_CSC_dl_for_check.scala 154:33:@120.4]
  reg [31:0] _RAND_16;
  reg [2:0] _T_872; // @[NV_NVDLA_CSC_dl_for_check.scala 155:29:@121.4]
  reg [31:0] _RAND_17;
  reg [2:0] _T_875; // @[NV_NVDLA_CSC_dl_for_check.scala 156:29:@122.4]
  reg [31:0] _RAND_18;
  reg [2:0] _T_881; // @[NV_NVDLA_CSC_dl_for_check.scala 158:29:@124.4]
  reg [31:0] _RAND_19;
  reg [2:0] _T_884; // @[NV_NVDLA_CSC_dl_for_check.scala 159:29:@125.4]
  reg [31:0] _RAND_20;
  reg [2:0] _T_887; // @[NV_NVDLA_CSC_dl_for_check.scala 160:29:@126.4]
  reg [31:0] _RAND_21;
  reg [2:0] _T_890; // @[NV_NVDLA_CSC_dl_for_check.scala 161:29:@127.4]
  reg [31:0] _RAND_22;
  reg [2:0] _T_896; // @[NV_NVDLA_CSC_dl_for_check.scala 163:29:@129.4]
  reg [31:0] _RAND_23;
  reg [2:0] _T_899; // @[NV_NVDLA_CSC_dl_for_check.scala 164:29:@130.4]
  reg [31:0] _RAND_24;
  reg [2:0] _T_905; // @[NV_NVDLA_CSC_dl_for_check.scala 166:30:@132.4]
  reg [31:0] _RAND_25;
  reg [2:0] _T_908; // @[NV_NVDLA_CSC_dl_for_check.scala 167:27:@133.4]
  reg [31:0] _RAND_26;
  reg [2:0] _T_911; // @[NV_NVDLA_CSC_dl_for_check.scala 168:27:@134.4]
  reg [31:0] _RAND_27;
  reg [3:0] _T_918; // @[NV_NVDLA_CSC_dl_for_check.scala 169:28:@136.4]
  reg [31:0] _RAND_28;
  reg [3:0] _T_925; // @[NV_NVDLA_CSC_dl_for_check.scala 170:28:@138.4]
  reg [31:0] _RAND_29;
  reg [4:0] _T_935; // @[NV_NVDLA_CSC_dl_for_check.scala 172:24:@141.4]
  reg [31:0] _RAND_30;
  reg [6:0] _T_942; // @[NV_NVDLA_CSC_dl_for_check.scala 173:27:@143.4]
  reg [31:0] _RAND_31;
  reg [6:0] _T_949; // @[NV_NVDLA_CSC_dl_for_check.scala 174:34:@145.4]
  reg [31:0] _RAND_32;
  reg [7:0] _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 175:26:@147.4]
  reg [31:0] _RAND_33;
  reg [6:0] _T_963; // @[NV_NVDLA_CSC_dl_for_check.scala 176:34:@149.4]
  reg [31:0] _RAND_34;
  reg [11:0] _T_970; // @[NV_NVDLA_CSC_dl_for_check.scala 177:30:@151.4]
  reg [31:0] _RAND_35;
  reg [5:0] _T_977; // @[NV_NVDLA_CSC_dl_for_check.scala 178:23:@153.4]
  reg [31:0] _RAND_36;
  reg [5:0] _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 179:23:@155.4]
  reg [31:0] _RAND_37;
  reg [15:0] _T_991; // @[NV_NVDLA_CSC_dl_for_check.scala 180:24:@157.4]
  reg [31:0] _RAND_38;
  reg [14:0] _T_998; // @[NV_NVDLA_CSC_dl_for_check.scala 181:26:@159.4]
  reg [31:0] _RAND_39;
  reg [14:0] _T_1005; // @[NV_NVDLA_CSC_dl_for_check.scala 182:30:@161.4]
  reg [31:0] _RAND_40;
  reg [14:0] _T_1012; // @[NV_NVDLA_CSC_dl_for_check.scala 183:30:@163.4]
  reg [31:0] _RAND_41;
  reg [13:0] _T_1019; // @[NV_NVDLA_CSC_dl_for_check.scala 185:26:@165.4]
  reg [31:0] _RAND_42;
  reg [14:0] _T_1026; // @[NV_NVDLA_CSC_dl_for_check.scala 186:27:@167.4]
  reg [31:0] _RAND_43;
  wire [33:0] _T_1041; // @[Bitwise.scala 72:12:@175.6]
  wire [5:0] _T_1043; // @[NV_NVDLA_CSC_dl_for_check.scala 193:38:@177.6]
  wire [4:0] _T_1044; // @[NV_NVDLA_CSC_dl_for_check.scala 193:38:@178.6]
  wire [13:0] _T_1046; // @[NV_NVDLA_CSC_dl_for_check.scala 194:48:@180.6]
  wire [6:0] _T_1052; // @[NV_NVDLA_CSC_dl_for_check.scala 197:93:@185.6]
  wire [10:0] _T_1053; // @[Cat.scala 30:58:@186.6]
  wire [14:0] _T_1057; // @[Cat.scala 30:58:@219.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [4:0] _GEN_2; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [13:0] _GEN_3; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [12:0] _GEN_4; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [12:0] _GEN_5; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [10:0] _GEN_6; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_7; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_8; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_10; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_11; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_12; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_13; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_15; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_19; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [2:0] _GEN_20; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [3:0] _GEN_21; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [5:0] _GEN_24; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [6:0] _GEN_26; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [6:0] _GEN_27; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [11:0] _GEN_30; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [5:0] _GEN_31; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [14:0] _GEN_34; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [14:0] _GEN_35; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [14:0] _GEN_36; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [13:0] _GEN_37; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [13:0] _GEN_39; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [12:0] _GEN_40; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  wire [11:0] _GEN_43; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  wire [11:0] _GEN_44; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  wire [14:0] _GEN_45; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  wire [14:0] _GEN_46; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  wire [14:0] _GEN_47; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  wire [13:0] _GEN_48; // @[NV_NVDLA_CSC_dl_for_check.scala 242:17:@239.4]
  wire [14:0] _GEN_49; // @[NV_NVDLA_CSC_dl_for_check.scala 242:17:@239.4]
  reg [14:0] _T_1079; // @[NV_NVDLA_CSC_dl_for_check.scala 265:59:@251.4]
  reg [31:0] _RAND_44;
  wire  _T_1159; // @[NV_NVDLA_CSC_dl_for_check.scala 306:37:@314.4]
  wire  _T_1160; // @[NV_NVDLA_CSC_dl_for_check.scala 306:23:@315.4]
  wire  _T_2244; // @[NV_NVDLA_CSC_dl_for_check.scala 896:32:@1229.4]
  reg  _T_2220; // @[NV_NVDLA_CSC_dl_for_check.scala 881:41:@1197.4]
  reg [31:0] _RAND_45;
  wire  _T_2245; // @[NV_NVDLA_CSC_dl_for_check.scala 896:36:@1230.4]
  wire  _T_2246; // @[NV_NVDLA_CSC_dl_for_check.scala 897:35:@1231.4]
  reg  _T_2214; // @[NV_NVDLA_CSC_dl_for_check.scala 881:41:@1195.4]
  reg [31:0] _RAND_46;
  wire  _T_2247; // @[NV_NVDLA_CSC_dl_for_check.scala 897:39:@1232.4]
  wire  _T_2248; // @[NV_NVDLA_CSC_dl_for_check.scala 896:57:@1233.4]
  wire  _T_2249; // @[NV_NVDLA_CSC_dl_for_check.scala 898:35:@1234.4]
  reg  _T_2211; // @[NV_NVDLA_CSC_dl_for_check.scala 881:41:@1194.4]
  reg [31:0] _RAND_47;
  wire  _T_2250; // @[NV_NVDLA_CSC_dl_for_check.scala 898:39:@1235.4]
  wire  _T_2251; // @[NV_NVDLA_CSC_dl_for_check.scala 897:60:@1236.4]
  wire  _T_2252; // @[NV_NVDLA_CSC_dl_for_check.scala 905:42:@1238.4]
  wire [26:0] _T_2256; // @[Bitwise.scala 72:12:@1240.4]
  reg [26:0] _T_2234; // @[NV_NVDLA_CSC_dl_for_check.scala 883:41:@1202.4]
  reg [31:0] _RAND_48;
  wire [26:0] _T_2257; // @[NV_NVDLA_CSC_dl_for_check.scala 905:47:@1241.4]
  wire  _T_2258; // @[NV_NVDLA_CSC_dl_for_check.scala 906:42:@1242.4]
  wire [26:0] _T_2262; // @[Bitwise.scala 72:12:@1244.4]
  reg [26:0] _T_2228; // @[NV_NVDLA_CSC_dl_for_check.scala 883:41:@1200.4]
  reg [31:0] _RAND_49;
  wire [26:0] _T_2263; // @[NV_NVDLA_CSC_dl_for_check.scala 906:47:@1245.4]
  wire [26:0] _T_2264; // @[NV_NVDLA_CSC_dl_for_check.scala 905:66:@1246.4]
  wire  _T_2265; // @[NV_NVDLA_CSC_dl_for_check.scala 907:42:@1247.4]
  wire [26:0] _T_2269; // @[Bitwise.scala 72:12:@1249.4]
  reg [26:0] _T_2225; // @[NV_NVDLA_CSC_dl_for_check.scala 883:41:@1199.4]
  reg [31:0] _RAND_50;
  wire [26:0] _T_2270; // @[NV_NVDLA_CSC_dl_for_check.scala 907:47:@1250.4]
  wire [26:0] _T_2271; // @[NV_NVDLA_CSC_dl_for_check.scala 906:66:@1251.4]
  wire  _T_2290; // @[NV_NVDLA_CSC_dl_for_check.scala 931:26:@1270.4]
  wire  _T_1157; // @[NV_NVDLA_CSC_dl_for_check.scala 303:29:@313.4]
  wire  _T_1162; // @[NV_NVDLA_CSC_dl_for_check.scala 306:66:@316.4]
  wire  _T_1163; // @[NV_NVDLA_CSC_dl_for_check.scala 306:53:@317.4]
  wire  _T_1164; // @[NV_NVDLA_CSC_dl_for_check.scala 306:42:@318.4]
  wire [13:0] _T_1165; // @[NV_NVDLA_CSC_dl_for_check.scala 307:28:@320.4]
  wire [14:0] _T_1166; // @[NV_NVDLA_CSC_dl_for_check.scala 308:29:@322.4]
  wire [14:0] _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 275:28:@262.4]
  wire [15:0] _T_1105; // @[NV_NVDLA_CSC_dl_for_check.scala 280:37:@269.4]
  wire [14:0] _T_1106; // @[NV_NVDLA_CSC_dl_for_check.scala 280:37:@270.4]
  wire [13:0] _T_1112; // @[Cat.scala 30:58:@272.4]
  wire [14:0] _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@273.4]
  wire [15:0] _T_1113; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@273.4]
  wire [15:0] _T_1114; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@274.4]
  wire [14:0] _T_1115; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@275.4]
  wire  _T_1122; // @[NV_NVDLA_CSC_dl_for_check.scala 282:45:@278.4]
  wire [14:0] _T_1124; // @[NV_NVDLA_CSC_dl_for_check.scala 283:83:@279.4]
  wire [14:0] _T_1125; // @[NV_NVDLA_CSC_dl_for_check.scala 283:25:@280.4]
  wire  _T_1151; // @[NV_NVDLA_CSC_dl_for_check.scala 294:13:@303.4]
  wire [14:0] _GEN_52; // @[NV_NVDLA_CSC_dl_for_check.scala 294:25:@304.4]
  reg  _T_1169; // @[NV_NVDLA_CSC_dl_for_check.scala 310:37:@324.4]
  reg [31:0] _RAND_51;
  reg [13:0] _T_1172; // @[Reg.scala 19:20:@327.4]
  reg [31:0] _RAND_52;
  wire [13:0] _GEN_54; // @[Reg.scala 20:19:@328.4]
  reg [14:0] _T_1175; // @[Reg.scala 19:20:@332.4]
  reg [31:0] _RAND_53;
  wire [14:0] _GEN_55; // @[Reg.scala 20:19:@333.4]
  reg  _T_1180; // @[NV_NVDLA_CSC_dl_for_check.scala 323:50:@338.4]
  reg [31:0] _RAND_54;
  reg  _T_1183; // @[NV_NVDLA_CSC_dl_for_check.scala 323:50:@339.4]
  reg [31:0] _RAND_55;
  reg  _T_1186; // @[NV_NVDLA_CSC_dl_for_check.scala 323:50:@340.4]
  reg [31:0] _RAND_56;
  reg  _T_1189; // @[NV_NVDLA_CSC_dl_for_check.scala 323:50:@341.4]
  reg [31:0] _RAND_57;
  reg  _T_1192; // @[NV_NVDLA_CSC_dl_for_check.scala 323:50:@342.4]
  reg [31:0] _RAND_58;
  reg  _T_1214; // @[NV_NVDLA_CSC_dl_for_check.scala 342:36:@372.4]
  reg [31:0] _RAND_59;
  reg  _T_1217; // @[NV_NVDLA_CSC_dl_for_check.scala 342:36:@373.4]
  reg [31:0] _RAND_60;
  reg  _T_1220; // @[NV_NVDLA_CSC_dl_for_check.scala 342:36:@374.4]
  reg [31:0] _RAND_61;
  reg  _T_1223; // @[NV_NVDLA_CSC_dl_for_check.scala 342:36:@375.4]
  reg [31:0] _RAND_62;
  reg [30:0] _T_1228; // @[NV_NVDLA_CSC_dl_for_check.scala 344:34:@377.4]
  reg [31:0] _RAND_63;
  reg [30:0] _T_1231; // @[NV_NVDLA_CSC_dl_for_check.scala 344:34:@378.4]
  reg [31:0] _RAND_64;
  reg [30:0] _T_1234; // @[NV_NVDLA_CSC_dl_for_check.scala 344:34:@379.4]
  reg [31:0] _RAND_65;
  reg [30:0] _T_1237; // @[NV_NVDLA_CSC_dl_for_check.scala 344:34:@380.4]
  reg [31:0] _RAND_66;
  wire [30:0] _T_1225; // @[NV_NVDLA_CSC_dl_for_check.scala 343:19:@376.4 NV_NVDLA_CSC_dl_for_check.scala 347:12:@382.4]
  wire [30:0] _GEN_61; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@384.4]
  wire [30:0] _GEN_62; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@388.4]
  wire [30:0] _GEN_63; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@392.4]
  wire [30:0] _GEN_64; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@396.4]
  wire  _T_1238; // @[NV_NVDLA_CSC_dl_for_check.scala 356:30:@399.4]
  wire  _T_1239; // @[NV_NVDLA_CSC_dl_for_check.scala 356:34:@400.4]
  wire  _T_1240; // @[NV_NVDLA_CSC_dl_for_check.scala 357:30:@401.4]
  wire  _T_1241; // @[NV_NVDLA_CSC_dl_for_check.scala 357:34:@402.4]
  wire  _T_1242; // @[NV_NVDLA_CSC_dl_for_check.scala 356:50:@403.4]
  wire  _T_1243; // @[NV_NVDLA_CSC_dl_for_check.scala 358:30:@404.4]
  wire  _T_1244; // @[NV_NVDLA_CSC_dl_for_check.scala 358:34:@405.4]
  wire  _T_1245; // @[NV_NVDLA_CSC_dl_for_check.scala 357:50:@406.4]
  wire  _T_1246; // @[NV_NVDLA_CSC_dl_for_check.scala 360:37:@407.4]
  wire [30:0] _T_1250; // @[Bitwise.scala 72:12:@409.4]
  wire [30:0] _T_1251; // @[NV_NVDLA_CSC_dl_for_check.scala 360:42:@410.4]
  wire  _T_1252; // @[NV_NVDLA_CSC_dl_for_check.scala 361:37:@411.4]
  wire [30:0] _T_1256; // @[Bitwise.scala 72:12:@413.4]
  wire [30:0] _T_1257; // @[NV_NVDLA_CSC_dl_for_check.scala 361:42:@414.4]
  wire [30:0] _T_1258; // @[NV_NVDLA_CSC_dl_for_check.scala 360:56:@415.4]
  wire  _T_1259; // @[NV_NVDLA_CSC_dl_for_check.scala 362:37:@416.4]
  wire [30:0] _T_1263; // @[Bitwise.scala 72:12:@418.4]
  wire [30:0] _T_1264; // @[NV_NVDLA_CSC_dl_for_check.scala 362:42:@419.4]
  wire [30:0] _T_1265; // @[NV_NVDLA_CSC_dl_for_check.scala 361:56:@420.4]
  wire [4:0] _T_1266; // @[NV_NVDLA_CSC_dl_for_check.scala 365:24:@421.4]
  wire [4:0] _T_1267; // @[NV_NVDLA_CSC_dl_for_check.scala 366:24:@422.4]
  wire [6:0] _T_1268; // @[NV_NVDLA_CSC_dl_for_check.scala 367:28:@423.4]
  wire [6:0] _T_1269; // @[NV_NVDLA_CSC_dl_for_check.scala 368:29:@424.4]
  wire [1:0] _T_1270; // @[NV_NVDLA_CSC_dl_for_check.scala 369:25:@425.4]
  wire  _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 370:25:@426.4]
  wire  _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 371:27:@427.4]
  wire  _T_1273; // @[NV_NVDLA_CSC_dl_for_check.scala 372:25:@428.4]
  wire  _T_1274; // @[NV_NVDLA_CSC_dl_for_check.scala 373:25:@429.4]
  wire  _T_1275; // @[NV_NVDLA_CSC_dl_for_check.scala 374:27:@430.4]
  reg [4:0] _T_1282; // @[NV_NVDLA_CSC_dl_for_check.scala 379:24:@433.4]
  reg [31:0] _RAND_67;
  wire [5:0] _T_1286; // @[NV_NVDLA_CSC_dl_for_check.scala 383:24:@434.4]
  wire [4:0] _T_1287; // @[NV_NVDLA_CSC_dl_for_check.scala 383:24:@435.4]
  wire  _T_1290; // @[NV_NVDLA_CSC_dl_for_check.scala 385:27:@439.4]
  wire [4:0] _T_1288; // @[NV_NVDLA_CSC_dl_for_check.scala 382:17:@436.4]
  wire [4:0] _T_1289; // @[NV_NVDLA_CSC_dl_for_check.scala 381:17:@437.4]
  reg [1:0] _T_1293; // @[NV_NVDLA_CSC_dl_for_check.scala 388:24:@441.4]
  reg [31:0] _RAND_68;
  wire [2:0] _T_1297; // @[NV_NVDLA_CSC_dl_for_check.scala 391:31:@443.4]
  wire [1:0] _T_1298; // @[NV_NVDLA_CSC_dl_for_check.scala 391:31:@444.4]
  wire [2:0] _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 392:32:@445.4]
  wire  _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 392:32:@445.4]
  wire  _T_1301; // @[NV_NVDLA_CSC_dl_for_check.scala 393:61:@447.4]
  reg [6:0] _T_1309; // @[NV_NVDLA_CSC_dl_for_check.scala 399:25:@455.4]
  reg [31:0] _RAND_69;
  wire  _T_1349; // @[NV_NVDLA_CSC_dl_for_check.scala 426:37:@484.4]
  wire  _T_1350; // @[NV_NVDLA_CSC_dl_for_check.scala 426:24:@485.4]
  wire  _T_1352; // @[NV_NVDLA_CSC_dl_for_check.scala 426:56:@486.4]
  wire  _T_1353; // @[NV_NVDLA_CSC_dl_for_check.scala 426:44:@487.4]
  wire  _T_1354; // @[NV_NVDLA_CSC_dl_for_check.scala 426:42:@488.4]
  wire  _T_1356; // @[NV_NVDLA_CSC_dl_for_check.scala 426:75:@489.4]
  wire  _T_1357; // @[NV_NVDLA_CSC_dl_for_check.scala 426:63:@490.4]
  wire  _T_1358; // @[NV_NVDLA_CSC_dl_for_check.scala 426:61:@491.4]
  reg  _T_1338; // @[NV_NVDLA_CSC_dl_for_check.scala 418:32:@477.4]
  reg [31:0] _RAND_70;
  wire  _T_1360; // @[NV_NVDLA_CSC_dl_for_check.scala 426:22:@492.4]
  wire  _T_1361; // @[NV_NVDLA_CSC_dl_for_check.scala 425:22:@493.4]
  wire  _T_1302; // @[NV_NVDLA_CSC_dl_for_check.scala 393:66:@448.4]
  wire  _T_1303; // @[NV_NVDLA_CSC_dl_for_check.scala 393:33:@449.4]
  wire  _T_1304; // @[NV_NVDLA_CSC_dl_for_check.scala 395:31:@451.6]
  wire [1:0] _T_1306; // @[NV_NVDLA_CSC_dl_for_check.scala 395:21:@452.6]
  wire [1:0] _GEN_65; // @[NV_NVDLA_CSC_dl_for_check.scala 394:23:@450.4]
  wire [7:0] _T_1315; // @[NV_NVDLA_CSC_dl_for_check.scala 403:33:@458.4]
  wire [6:0] _T_1316; // @[NV_NVDLA_CSC_dl_for_check.scala 403:33:@459.4]
  wire  _T_1317; // @[NV_NVDLA_CSC_dl_for_check.scala 404:51:@460.4]
  wire  _T_1318; // @[NV_NVDLA_CSC_dl_for_check.scala 404:33:@461.4]
  wire  _T_1319; // @[NV_NVDLA_CSC_dl_for_check.scala 405:34:@463.4]
  wire  _T_1320; // @[NV_NVDLA_CSC_dl_for_check.scala 406:52:@465.4]
  wire  _T_1321; // @[NV_NVDLA_CSC_dl_for_check.scala 406:34:@466.4]
  wire  _T_1323; // @[NV_NVDLA_CSC_dl_for_check.scala 410:41:@468.6]
  wire  _T_1324; // @[NV_NVDLA_CSC_dl_for_check.scala 410:39:@469.6]
  wire [6:0] _T_1327; // @[NV_NVDLA_CSC_dl_for_check.scala 411:22:@470.6]
  wire [6:0] _T_1328; // @[NV_NVDLA_CSC_dl_for_check.scala 410:22:@471.6]
  wire [6:0] _T_1329; // @[NV_NVDLA_CSC_dl_for_check.scala 409:22:@472.6]
  wire [6:0] _GEN_66; // @[NV_NVDLA_CSC_dl_for_check.scala 408:24:@467.4]
  reg  _T_1332; // @[NV_NVDLA_CSC_dl_for_check.scala 416:35:@475.4]
  reg [31:0] _RAND_71;
  reg  _T_1335; // @[NV_NVDLA_CSC_dl_for_check.scala 417:32:@476.4]
  reg [31:0] _RAND_72;
  wire  _T_1346; // @[NV_NVDLA_CSC_dl_for_check.scala 424:27:@482.4]
  wire  _T_1341; // @[NV_NVDLA_CSC_dl_for_check.scala 421:49:@479.4]
  wire  _T_1344; // @[NV_NVDLA_CSC_dl_for_check.scala 422:32:@480.4]
  wire  _T_1345; // @[NV_NVDLA_CSC_dl_for_check.scala 421:33:@481.4]
  reg [7:0] _T_1364; // @[NV_NVDLA_CSC_dl_for_check.scala 434:31:@498.4]
  reg [31:0] _RAND_73;
  wire [7:0] _T_1366; // @[Cat.scala 30:58:@499.4]
  wire [7:0] _GEN_67; // @[NV_NVDLA_CSC_dl_for_check.scala 436:21:@500.4]
  reg [12:0] _T_1369; // @[NV_NVDLA_CSC_dl_for_check.scala 442:28:@503.4]
  reg [31:0] _RAND_74;
  reg [12:0] _T_1372; // @[NV_NVDLA_CSC_dl_for_check.scala 443:28:@504.4]
  reg [31:0] _RAND_75;
  wire [12:0] _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 446:39:@505.4]
  wire [13:0] _T_1373; // @[NV_NVDLA_CSC_dl_for_check.scala 446:39:@505.4]
  wire [12:0] _T_1374; // @[NV_NVDLA_CSC_dl_for_check.scala 446:39:@506.4]
  wire  _T_1375; // @[NV_NVDLA_CSC_dl_for_check.scala 447:29:@507.4]
  wire  _T_1376; // @[NV_NVDLA_CSC_dl_for_check.scala 447:61:@508.4]
  wire  _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 447:44:@509.4]
  wire  _T_1380; // @[NV_NVDLA_CSC_dl_for_check.scala 450:43:@512.4]
  wire  _T_1381; // @[NV_NVDLA_CSC_dl_for_check.scala 450:41:@513.4]
  wire [12:0] _T_1382; // @[NV_NVDLA_CSC_dl_for_check.scala 451:26:@514.4]
  wire [12:0] _T_1383; // @[NV_NVDLA_CSC_dl_for_check.scala 450:26:@515.4]
  wire [12:0] _T_1384; // @[NV_NVDLA_CSC_dl_for_check.scala 449:26:@516.4]
  wire  _T_1386; // @[NV_NVDLA_CSC_dl_for_check.scala 452:70:@518.4]
  wire  _T_1387; // @[NV_NVDLA_CSC_dl_for_check.scala 452:37:@519.4]
  wire  _T_1388; // @[NV_NVDLA_CSC_dl_for_check.scala 453:55:@520.4]
  wire  _T_1389; // @[NV_NVDLA_CSC_dl_for_check.scala 453:71:@521.4]
  wire  _T_1390; // @[NV_NVDLA_CSC_dl_for_check.scala 453:37:@522.4]
  wire [12:0] _GEN_68; // @[NV_NVDLA_CSC_dl_for_check.scala 455:27:@523.4]
  wire [12:0] _GEN_69; // @[NV_NVDLA_CSC_dl_for_check.scala 458:27:@526.4]
  reg [10:0] _T_1393; // @[NV_NVDLA_CSC_dl_for_check.scala 463:27:@529.4]
  reg [31:0] _RAND_76;
  wire  _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 465:37:@530.4]
  wire  _T_1396; // @[NV_NVDLA_CSC_dl_for_check.scala 466:70:@532.4]
  wire  _T_1397; // @[NV_NVDLA_CSC_dl_for_check.scala 466:36:@533.4]
  wire [11:0] _T_1401; // @[NV_NVDLA_CSC_dl_for_check.scala 471:34:@535.6]
  wire [10:0] _T_1402; // @[NV_NVDLA_CSC_dl_for_check.scala 471:34:@536.6]
  wire [10:0] _T_1403; // @[NV_NVDLA_CSC_dl_for_check.scala 470:24:@537.6]
  wire [10:0] _T_1404; // @[NV_NVDLA_CSC_dl_for_check.scala 469:24:@538.6]
  wire [10:0] _GEN_70; // @[NV_NVDLA_CSC_dl_for_check.scala 468:26:@534.4]
  reg [13:0] _T_1407; // @[NV_NVDLA_CSC_dl_for_check.scala 475:27:@541.4]
  reg [31:0] _RAND_77;
  reg [13:0] _T_1410; // @[NV_NVDLA_CSC_dl_for_check.scala 476:27:@542.4]
  reg [31:0] _RAND_78;
  reg [15:0] _T_1413; // @[NV_NVDLA_CSC_dl_for_check.scala 477:26:@543.4]
  reg [31:0] _RAND_79;
  reg [15:0] _T_1416; // @[NV_NVDLA_CSC_dl_for_check.scala 478:26:@544.4]
  reg [31:0] _RAND_80;
  reg [15:0] _T_1419; // @[NV_NVDLA_CSC_dl_for_check.scala 479:29:@545.4]
  reg [31:0] _RAND_81;
  reg [12:0] _T_1422; // @[NV_NVDLA_CSC_dl_for_check.scala 480:29:@546.4]
  reg [31:0] _RAND_82;
  reg  _T_1427; // @[NV_NVDLA_CSC_dl_for_check.scala 482:33:@548.4]
  reg [31:0] _RAND_83;
  reg  _T_1430; // @[NV_NVDLA_CSC_dl_for_check.scala 483:35:@549.4]
  reg [31:0] _RAND_84;
  wire [12:0] _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 486:41:@550.4]
  wire [13:0] _T_1433; // @[NV_NVDLA_CSC_dl_for_check.scala 486:41:@550.4]
  wire [13:0] _T_1434; // @[NV_NVDLA_CSC_dl_for_check.scala 486:41:@551.4]
  wire [13:0] _T_1435; // @[NV_NVDLA_CSC_dl_for_check.scala 485:26:@552.4]
  wire [13:0] _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@553.4]
  wire [14:0] _T_1436; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@553.4]
  wire [13:0] _T_1437; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@554.4]
  wire [13:0] _T_1440; // @[NV_NVDLA_CSC_dl_for_check.scala 492:25:@557.4]
  wire [13:0] _T_1441; // @[NV_NVDLA_CSC_dl_for_check.scala 491:25:@558.4]
  wire [13:0] _T_1442; // @[NV_NVDLA_CSC_dl_for_check.scala 490:25:@559.4]
  wire [5:0] _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 494:35:@560.4]
  wire [10:0] _T_1443; // @[NV_NVDLA_CSC_dl_for_check.scala 494:35:@560.4]
  wire [13:0] _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@561.4]
  wire [14:0] _T_1444; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@561.4]
  wire [13:0] _T_1445; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@562.4]
  wire  _T_1448; // @[NV_NVDLA_CSC_dl_for_check.scala 496:96:@565.4]
  wire  _T_1449; // @[NV_NVDLA_CSC_dl_for_check.scala 496:86:@566.4]
  wire  _T_1450; // @[NV_NVDLA_CSC_dl_for_check.scala 496:84:@567.4]
  wire  _T_1451; // @[NV_NVDLA_CSC_dl_for_check.scala 496:36:@568.4]
  wire  _T_1454; // @[NV_NVDLA_CSC_dl_for_check.scala 497:99:@571.4]
  wire  _T_1455; // @[NV_NVDLA_CSC_dl_for_check.scala 497:89:@572.4]
  wire  _T_1456; // @[NV_NVDLA_CSC_dl_for_check.scala 497:87:@573.4]
  wire  _T_1457; // @[NV_NVDLA_CSC_dl_for_check.scala 497:36:@574.4]
  wire [7:0] _T_1459; // @[NV_NVDLA_CSC_dl_for_check.scala 500:26:@575.4]
  wire  _T_1462; // @[NV_NVDLA_CSC_dl_for_check.scala 502:79:@577.4]
  wire [7:0] _T_1466; // @[NV_NVDLA_CSC_dl_for_check.scala 503:74:@580.4]
  wire [6:0] _T_1467; // @[NV_NVDLA_CSC_dl_for_check.scala 503:74:@581.4]
  wire [6:0] _T_1468; // @[NV_NVDLA_CSC_dl_for_check.scala 502:27:@582.4]
  wire  _T_1469; // @[NV_NVDLA_CSC_dl_for_check.scala 504:37:@583.4]
  wire  _T_1471; // @[NV_NVDLA_CSC_dl_for_check.scala 505:35:@584.4]
  wire [13:0] _T_1473; // @[NV_NVDLA_CSC_dl_for_check.scala 505:66:@585.4]
  wire [12:0] _T_1474; // @[NV_NVDLA_CSC_dl_for_check.scala 505:66:@586.4]
  wire [12:0] _T_1475; // @[NV_NVDLA_CSC_dl_for_check.scala 505:22:@587.4]
  wire [12:0] _T_1476; // @[NV_NVDLA_CSC_dl_for_check.scala 504:22:@588.4]
  wire [12:0] _GEN_688; // @[NV_NVDLA_CSC_dl_for_check.scala 507:44:@590.4]
  wire  _T_1477; // @[NV_NVDLA_CSC_dl_for_check.scala 507:44:@590.4]
  wire  _T_1478; // @[NV_NVDLA_CSC_dl_for_check.scala 511:39:@591.4]
  wire  _T_1479; // @[NV_NVDLA_CSC_dl_for_check.scala 511:54:@592.4]
  wire  _T_1480; // @[NV_NVDLA_CSC_dl_for_check.scala 511:71:@593.4]
  wire  _T_1483; // @[NV_NVDLA_CSC_dl_for_check.scala 512:73:@596.4]
  wire  _T_1484; // @[NV_NVDLA_CSC_dl_for_check.scala 512:71:@597.4]
  wire [15:0] _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 512:99:@598.4]
  wire [16:0] _T_1485; // @[NV_NVDLA_CSC_dl_for_check.scala 512:99:@598.4]
  wire [15:0] _T_1486; // @[NV_NVDLA_CSC_dl_for_check.scala 512:99:@599.4]
  wire  _T_1488; // @[NV_NVDLA_CSC_dl_for_check.scala 513:54:@601.4]
  wire [15:0] _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 513:90:@602.4]
  wire [16:0] _T_1489; // @[NV_NVDLA_CSC_dl_for_check.scala 513:90:@602.4]
  wire [15:0] _T_1490; // @[NV_NVDLA_CSC_dl_for_check.scala 513:90:@603.4]
  wire  _T_1492; // @[NV_NVDLA_CSC_dl_for_check.scala 514:56:@605.4]
  wire  _T_1493; // @[NV_NVDLA_CSC_dl_for_check.scala 514:54:@606.4]
  wire [16:0] _T_1495; // @[NV_NVDLA_CSC_dl_for_check.scala 514:91:@607.4]
  wire [15:0] _T_1496; // @[NV_NVDLA_CSC_dl_for_check.scala 514:91:@608.4]
  wire  _T_1497; // @[NV_NVDLA_CSC_dl_for_check.scala 515:41:@609.4]
  wire  _T_1498; // @[NV_NVDLA_CSC_dl_for_check.scala 515:39:@610.4]
  wire [15:0] _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 515:81:@611.4]
  wire [16:0] _T_1499; // @[NV_NVDLA_CSC_dl_for_check.scala 515:81:@611.4]
  wire [15:0] _T_1500; // @[NV_NVDLA_CSC_dl_for_check.scala 515:81:@612.4]
  wire [15:0] _T_1501; // @[NV_NVDLA_CSC_dl_for_check.scala 515:24:@613.4]
  wire [15:0] _T_1502; // @[NV_NVDLA_CSC_dl_for_check.scala 514:24:@614.4]
  wire [15:0] _T_1503; // @[NV_NVDLA_CSC_dl_for_check.scala 513:24:@615.4]
  wire [15:0] _T_1504; // @[NV_NVDLA_CSC_dl_for_check.scala 512:24:@616.4]
  wire [15:0] _T_1505; // @[NV_NVDLA_CSC_dl_for_check.scala 511:24:@617.4]
  wire [15:0] _T_1506; // @[NV_NVDLA_CSC_dl_for_check.scala 510:24:@618.4]
  wire [9:0] _T_1512; // @[NV_NVDLA_CSC_dl_for_check.scala 517:68:@620.4]
  wire [14:0] _T_1513; // @[Cat.scala 30:58:@621.4]
  wire  _T_1524; // @[NV_NVDLA_CSC_dl_for_check.scala 520:68:@632.4]
  wire  _T_1525; // @[NV_NVDLA_CSC_dl_for_check.scala 520:57:@633.4]
  wire  _T_1526; // @[NV_NVDLA_CSC_dl_for_check.scala 520:72:@634.4]
  wire  _T_1527; // @[NV_NVDLA_CSC_dl_for_check.scala 520:88:@635.4]
  wire  _T_1528; // @[NV_NVDLA_CSC_dl_for_check.scala 520:103:@636.4]
  wire  _T_1529; // @[NV_NVDLA_CSC_dl_for_check.scala 520:39:@637.4]
  wire  _T_1531; // @[NV_NVDLA_CSC_dl_for_check.scala 522:42:@639.4]
  wire  _T_1534; // @[NV_NVDLA_CSC_dl_for_check.scala 522:74:@640.4]
  wire  _T_1535; // @[NV_NVDLA_CSC_dl_for_check.scala 522:28:@641.4]
  wire  _T_1537; // @[NV_NVDLA_CSC_dl_for_check.scala 523:36:@643.4]
  wire  _T_1538; // @[NV_NVDLA_CSC_dl_for_check.scala 523:72:@644.4]
  wire  _T_1539; // @[NV_NVDLA_CSC_dl_for_check.scala 523:51:@645.4]
  wire [13:0] _GEN_71; // @[NV_NVDLA_CSC_dl_for_check.scala 525:26:@646.4]
  wire [15:0] _GEN_72; // @[NV_NVDLA_CSC_dl_for_check.scala 525:26:@646.4]
  wire [13:0] _GEN_73; // @[NV_NVDLA_CSC_dl_for_check.scala 529:26:@650.4]
  wire [15:0] _GEN_74; // @[NV_NVDLA_CSC_dl_for_check.scala 529:26:@650.4]
  wire [15:0] _GEN_75; // @[NV_NVDLA_CSC_dl_for_check.scala 533:26:@654.4]
  reg [13:0] _T_1542; // @[NV_NVDLA_CSC_dl_for_check.scala 539:27:@657.4]
  reg [31:0] _RAND_85;
  reg [13:0] _T_1545; // @[NV_NVDLA_CSC_dl_for_check.scala 540:27:@658.4]
  reg [31:0] _RAND_86;
  wire [13:0] _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@659.4]
  wire [14:0] _T_1547; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@659.4]
  wire [14:0] _T_1548; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@660.4]
  wire [13:0] _T_1549; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@661.4]
  wire [13:0] _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 543:37:@662.4]
  wire [14:0] _T_1550; // @[NV_NVDLA_CSC_dl_for_check.scala 543:37:@662.4]
  wire [13:0] _T_1551; // @[NV_NVDLA_CSC_dl_for_check.scala 543:37:@663.4]
  wire  _T_1552; // @[NV_NVDLA_CSC_dl_for_check.scala 544:52:@664.4]
  wire  _T_1553; // @[NV_NVDLA_CSC_dl_for_check.scala 544:35:@665.4]
  wire [13:0] _T_1556; // @[NV_NVDLA_CSC_dl_for_check.scala 546:25:@668.4]
  wire [13:0] _T_1557; // @[NV_NVDLA_CSC_dl_for_check.scala 545:25:@669.4]
  wire [13:0] _T_1558; // @[NV_NVDLA_CSC_dl_for_check.scala 544:25:@670.4]
  wire  _T_1561; // @[NV_NVDLA_CSC_dl_for_check.scala 547:91:@673.4]
  wire  _T_1562; // @[NV_NVDLA_CSC_dl_for_check.scala 547:54:@674.4]
  wire  _T_1563; // @[NV_NVDLA_CSC_dl_for_check.scala 547:36:@675.4]
  wire [5:0] _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 549:35:@679.4]
  wire [10:0] _T_1567; // @[NV_NVDLA_CSC_dl_for_check.scala 549:35:@679.4]
  wire [13:0] _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 550:33:@680.4]
  wire [14:0] _T_1568; // @[NV_NVDLA_CSC_dl_for_check.scala 550:33:@680.4]
  wire [13:0] _T_1569; // @[NV_NVDLA_CSC_dl_for_check.scala 550:33:@681.4]
  wire [13:0] _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 550:51:@682.4]
  wire [14:0] _T_1570; // @[NV_NVDLA_CSC_dl_for_check.scala 550:51:@682.4]
  wire [13:0] _T_1571; // @[NV_NVDLA_CSC_dl_for_check.scala 550:51:@683.4]
  wire [13:0] _GEN_76; // @[NV_NVDLA_CSC_dl_for_check.scala 552:26:@684.4]
  wire [13:0] _GEN_77; // @[NV_NVDLA_CSC_dl_for_check.scala 553:26:@687.4]
  wire  _T_1572; // @[NV_NVDLA_CSC_dl_for_check.scala 556:39:@690.4]
  wire [13:0] _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 556:59:@691.4]
  wire  _T_1573; // @[NV_NVDLA_CSC_dl_for_check.scala 556:59:@691.4]
  wire  _T_1574; // @[NV_NVDLA_CSC_dl_for_check.scala 556:44:@692.4]
  wire  _T_1575; // @[NV_NVDLA_CSC_dl_for_check.scala 556:92:@693.4]
  wire  _T_1576; // @[NV_NVDLA_CSC_dl_for_check.scala 556:78:@694.4]
  wire [13:0] _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 556:112:@695.4]
  wire  _T_1577; // @[NV_NVDLA_CSC_dl_for_check.scala 556:112:@695.4]
  wire  _T_1578; // @[NV_NVDLA_CSC_dl_for_check.scala 556:97:@696.4]
  wire  _T_1591; // @[NV_NVDLA_CSC_dl_for_check.scala 559:42:@706.4]
  wire  _T_1701; // @[NV_NVDLA_CSC_dl_for_check.scala 644:33:@792.4]
  wire  _T_1702; // @[NV_NVDLA_CSC_dl_for_check.scala 645:24:@793.4]
  wire [12:0] _T_1704; // @[NV_NVDLA_CSC_dl_for_check.scala 645:77:@794.4]
  wire [14:0] _T_1705; // @[Cat.scala 30:58:@795.4]
  wire  _T_1707; // @[NV_NVDLA_CSC_dl_for_check.scala 646:38:@796.4]
  wire [11:0] _T_1712; // @[NV_NVDLA_CSC_dl_for_check.scala 647:54:@799.4]
  wire [14:0] _T_1713; // @[Cat.scala 30:58:@800.4]
  wire [14:0] _T_1714; // @[NV_NVDLA_CSC_dl_for_check.scala 646:23:@801.4]
  wire [14:0] _T_1715; // @[NV_NVDLA_CSC_dl_for_check.scala 645:23:@802.4]
  wire [14:0] _T_1716; // @[NV_NVDLA_CSC_dl_for_check.scala 644:23:@803.4]
  wire [13:0] _T_1717; // @[NV_NVDLA_CSC_dl_for_check.scala 656:24:@805.4]
  wire [11:0] _T_1594; // @[NV_NVDLA_CSC_dl_for_check.scala 563:32:@708.4]
  wire [14:0] _GEN_700; // @[NV_NVDLA_CSC_dl_for_check.scala 563:40:@709.4]
  wire  _T_1595; // @[NV_NVDLA_CSC_dl_for_check.scala 563:40:@709.4]
  wire  _T_1596; // @[NV_NVDLA_CSC_dl_for_check.scala 564:34:@710.4]
  wire  _T_1597; // @[NV_NVDLA_CSC_dl_for_check.scala 564:24:@711.4]
  wire  _T_1598; // @[NV_NVDLA_CSC_dl_for_check.scala 565:29:@712.4]
  wire  _T_1599; // @[NV_NVDLA_CSC_dl_for_check.scala 565:33:@713.4]
  wire  _T_1600; // @[NV_NVDLA_CSC_dl_for_check.scala 566:39:@714.4]
  wire  _T_1601; // @[NV_NVDLA_CSC_dl_for_check.scala 566:37:@715.4]
  wire  _T_1602; // @[NV_NVDLA_CSC_dl_for_check.scala 566:56:@716.4]
  wire  _T_1603; // @[NV_NVDLA_CSC_dl_for_check.scala 566:54:@717.4]
  wire  _T_1604; // @[NV_NVDLA_CSC_dl_for_check.scala 569:37:@718.4]
  wire  _T_1605; // @[NV_NVDLA_CSC_dl_for_check.scala 569:27:@719.4]
  wire  _T_1606; // @[NV_NVDLA_CSC_dl_for_check.scala 569:54:@720.4]
  wire  _T_1607; // @[NV_NVDLA_CSC_dl_for_check.scala 569:26:@721.4]
  wire [1:0] _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 570:35:@722.4]
  wire  _T_1610; // @[NV_NVDLA_CSC_dl_for_check.scala 571:55:@723.4]
  wire  _T_1611; // @[NV_NVDLA_CSC_dl_for_check.scala 571:42:@724.4]
  wire  _T_1612; // @[NV_NVDLA_CSC_dl_for_check.scala 574:42:@726.4]
  wire [8:0] _T_1616; // @[Cat.scala 30:58:@730.4]
  reg  _T_1619; // @[NV_NVDLA_CSC_dl_for_check.scala 581:31:@731.4]
  reg [31:0] _RAND_87;
  reg [1:0] _T_1622; // @[NV_NVDLA_CSC_dl_for_check.scala 582:31:@732.4]
  reg [31:0] _RAND_88;
  reg [1:0] _T_1625; // @[NV_NVDLA_CSC_dl_for_check.scala 583:31:@733.4]
  reg [31:0] _RAND_89;
  reg  _T_1628; // @[NV_NVDLA_CSC_dl_for_check.scala 584:31:@734.4]
  reg [31:0] _RAND_90;
  reg  _T_1631; // @[NV_NVDLA_CSC_dl_for_check.scala 585:32:@735.4]
  reg [31:0] _RAND_91;
  reg  _T_1634; // @[NV_NVDLA_CSC_dl_for_check.scala 586:31:@736.4]
  reg [31:0] _RAND_92;
  reg [1:0] _T_1637; // @[NV_NVDLA_CSC_dl_for_check.scala 587:35:@737.4]
  reg [31:0] _RAND_93;
  reg  _T_1640; // @[NV_NVDLA_CSC_dl_for_check.scala 588:34:@738.4]
  reg [31:0] _RAND_94;
  reg [8:0] _T_1643; // @[NV_NVDLA_CSC_dl_for_check.scala 589:30:@739.4]
  reg [31:0] _RAND_95;
  reg  _T_1646; // @[NV_NVDLA_CSC_dl_for_check.scala 590:29:@740.4]
  reg [31:0] _RAND_96;
  wire  _T_1647; // @[NV_NVDLA_CSC_dl_for_check.scala 601:38:@750.6]
  wire  _T_1648; // @[NV_NVDLA_CSC_dl_for_check.scala 601:56:@751.6]
  wire [1:0] _GEN_78; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire [1:0] _GEN_79; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_80; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_81; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_82; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire [1:0] _GEN_83; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire [8:0] _GEN_84; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_85; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_86; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_87; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  wire  _GEN_88; // @[NV_NVDLA_CSC_dl_for_check.scala 605:26:@756.4]
  reg [12:0] _T_1651; // @[NV_NVDLA_CSC_dl_for_check.scala 613:21:@759.4]
  reg [31:0] _RAND_97;
  reg [12:0] _T_1654; // @[NV_NVDLA_CSC_dl_for_check.scala 614:24:@760.4]
  reg [31:0] _RAND_98;
  reg [12:0] _T_1657; // @[NV_NVDLA_CSC_dl_for_check.scala 615:26:@761.4]
  reg [31:0] _RAND_99;
  reg [12:0] _T_1660; // @[NV_NVDLA_CSC_dl_for_check.scala 616:26:@762.4]
  reg [31:0] _RAND_100;
  reg [12:0] _T_1663; // @[NV_NVDLA_CSC_dl_for_check.scala 617:26:@763.4]
  reg [31:0] _RAND_101;
  reg [12:0] _T_1666; // @[NV_NVDLA_CSC_dl_for_check.scala 618:26:@764.4]
  reg [31:0] _RAND_102;
  reg [12:0] _T_1669; // @[NV_NVDLA_CSC_dl_for_check.scala 619:24:@765.4]
  reg [31:0] _RAND_103;
  wire  _T_1670; // @[NV_NVDLA_CSC_dl_for_check.scala 622:32:@766.4]
  wire  _T_1671; // @[NV_NVDLA_CSC_dl_for_check.scala 622:22:@767.4]
  wire [11:0] _T_1672; // @[NV_NVDLA_CSC_dl_for_check.scala 622:49:@768.4]
  wire [11:0] _T_1674; // @[NV_NVDLA_CSC_dl_for_check.scala 622:21:@769.4]
  wire  _T_1676; // @[NV_NVDLA_CSC_dl_for_check.scala 624:34:@770.4]
  wire [12:0] _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 624:64:@771.4]
  wire [13:0] _T_1678; // @[NV_NVDLA_CSC_dl_for_check.scala 624:64:@771.4]
  wire [12:0] _T_1679; // @[NV_NVDLA_CSC_dl_for_check.scala 624:64:@772.4]
  wire [12:0] _T_1680; // @[NV_NVDLA_CSC_dl_for_check.scala 624:19:@773.4]
  wire [12:0] _T_1681; // @[NV_NVDLA_CSC_dl_for_check.scala 623:19:@774.4]
  wire  _T_1685; // @[NV_NVDLA_CSC_dl_for_check.scala 626:31:@778.4]
  wire [13:0] _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 629:32:@779.4]
  wire [25:0] _T_1686; // @[NV_NVDLA_CSC_dl_for_check.scala 629:32:@779.4]
  wire [12:0] _T_1687; // @[NV_NVDLA_CSC_dl_for_check.scala 629:50:@780.4]
  wire [11:0] _GEN_703; // @[NV_NVDLA_CSC_dl_for_check.scala 630:31:@781.4]
  wire [16:0] _T_1688; // @[NV_NVDLA_CSC_dl_for_check.scala 630:31:@781.4]
  wire [12:0] _T_1689; // @[NV_NVDLA_CSC_dl_for_check.scala 630:49:@782.4]
  wire [14:0] _GEN_704; // @[NV_NVDLA_CSC_dl_for_check.scala 631:29:@783.4]
  wire [19:0] _T_1690; // @[NV_NVDLA_CSC_dl_for_check.scala 631:29:@783.4]
  wire [12:0] _T_1691; // @[NV_NVDLA_CSC_dl_for_check.scala 631:47:@784.4]
  wire [14:0] _GEN_705; // @[NV_NVDLA_CSC_dl_for_check.scala 632:47:@785.4]
  wire [16:0] _T_1693; // @[NV_NVDLA_CSC_dl_for_check.scala 632:47:@785.4]
  wire [16:0] _T_1694; // @[NV_NVDLA_CSC_dl_for_check.scala 632:21:@786.4]
  wire [12:0] _T_1695; // @[NV_NVDLA_CSC_dl_for_check.scala 632:65:@787.4]
  wire  _T_1696; // @[NV_NVDLA_CSC_dl_for_check.scala 633:45:@788.4]
  wire  _T_1697; // @[NV_NVDLA_CSC_dl_for_check.scala 633:34:@789.4]
  wire [1:0] _T_1698; // @[Cat.scala 30:58:@790.4]
  wire [12:0] _GEN_89; // @[NV_NVDLA_CSC_dl_for_check.scala 660:20:@807.4]
  wire [12:0] _GEN_90; // @[NV_NVDLA_CSC_dl_for_check.scala 663:23:@810.4]
  wire  _T_1718; // @[NV_NVDLA_CSC_dl_for_check.scala 666:19:@813.4]
  wire [12:0] _GEN_91; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@814.4]
  wire [12:0] _GEN_92; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@814.4]
  wire [12:0] _GEN_93; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@814.4]
  wire  _T_1719; // @[NV_NVDLA_CSC_dl_for_check.scala 671:19:@819.4]
  wire [12:0] _GEN_94; // @[NV_NVDLA_CSC_dl_for_check.scala 671:23:@820.4]
  wire [13:0] _GEN_95; // @[NV_NVDLA_CSC_dl_for_check.scala 674:20:@823.4]
  reg [12:0] _T_1762_0; // @[NV_NVDLA_CSC_dl_for_check.scala 682:33:@835.4]
  reg [31:0] _RAND_104;
  reg [12:0] _T_1762_1; // @[NV_NVDLA_CSC_dl_for_check.scala 682:33:@835.4]
  reg [31:0] _RAND_105;
  reg [12:0] _T_1762_2; // @[NV_NVDLA_CSC_dl_for_check.scala 682:33:@835.4]
  reg [31:0] _RAND_106;
  reg [12:0] _T_1762_3; // @[NV_NVDLA_CSC_dl_for_check.scala 682:33:@835.4]
  reg [31:0] _RAND_107;
  reg  _T_1781; // @[NV_NVDLA_CSC_dl_for_check.scala 683:35:@836.4]
  reg [31:0] _RAND_108;
  reg [14:0] _T_1788; // @[NV_NVDLA_CSC_dl_for_check.scala 684:37:@838.4]
  reg [31:0] _RAND_109;
  reg  _T_1791; // @[NV_NVDLA_CSC_dl_for_check.scala 685:32:@839.4]
  reg [31:0] _RAND_110;
  reg [1:0] _T_1797; // @[NV_NVDLA_CSC_dl_for_check.scala 687:33:@841.4]
  reg [31:0] _RAND_111;
  reg [1:0] _T_1800; // @[NV_NVDLA_CSC_dl_for_check.scala 688:33:@842.4]
  reg [31:0] _RAND_112;
  reg  _T_1803; // @[NV_NVDLA_CSC_dl_for_check.scala 689:33:@843.4]
  reg [31:0] _RAND_113;
  reg  _T_1806; // @[NV_NVDLA_CSC_dl_for_check.scala 690:34:@844.4]
  reg [31:0] _RAND_114;
  reg [7:0] _T_1809; // @[NV_NVDLA_CSC_dl_for_check.scala 691:33:@845.4]
  reg [31:0] _RAND_115;
  reg  _T_1812; // @[NV_NVDLA_CSC_dl_for_check.scala 692:33:@846.4]
  reg [31:0] _RAND_116;
  reg [1:0] _T_1815; // @[NV_NVDLA_CSC_dl_for_check.scala 693:37:@847.4]
  reg [31:0] _RAND_117;
  reg  _T_1818; // @[NV_NVDLA_CSC_dl_for_check.scala 694:36:@848.4]
  reg [31:0] _RAND_118;
  reg  _T_1821; // @[NV_NVDLA_CSC_dl_for_check.scala 695:31:@849.4]
  reg [31:0] _RAND_119;
  reg [8:0] _T_1824; // @[NV_NVDLA_CSC_dl_for_check.scala 696:32:@850.4]
  reg [31:0] _RAND_120;
  wire [13:0] _T_1825; // @[NV_NVDLA_CSC_dl_for_check.scala 698:29:@851.4]
  wire [12:0] _T_1826; // @[NV_NVDLA_CSC_dl_for_check.scala 698:29:@852.4]
  wire [13:0] _T_1827; // @[NV_NVDLA_CSC_dl_for_check.scala 698:43:@853.4]
  wire [12:0] _T_1828; // @[NV_NVDLA_CSC_dl_for_check.scala 698:43:@854.4]
  wire [13:0] _T_1829; // @[NV_NVDLA_CSC_dl_for_check.scala 698:57:@855.4]
  wire [12:0] _T_1830; // @[NV_NVDLA_CSC_dl_for_check.scala 698:57:@856.4]
  wire [14:0] _GEN_706; // @[NV_NVDLA_CSC_dl_for_check.scala 699:40:@857.4]
  wire [15:0] _T_1831; // @[NV_NVDLA_CSC_dl_for_check.scala 699:40:@857.4]
  wire [14:0] _T_1832; // @[NV_NVDLA_CSC_dl_for_check.scala 699:40:@858.4]
  wire [14:0] _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 699:52:@859.4]
  wire [15:0] _T_1833; // @[NV_NVDLA_CSC_dl_for_check.scala 699:52:@859.4]
  wire [14:0] _T_1834; // @[NV_NVDLA_CSC_dl_for_check.scala 699:52:@860.4]
  wire [14:0] _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 699:64:@861.4]
  wire [15:0] _T_1835; // @[NV_NVDLA_CSC_dl_for_check.scala 699:64:@861.4]
  wire [14:0] _T_1836; // @[NV_NVDLA_CSC_dl_for_check.scala 699:64:@862.4]
  wire  _T_1843; // @[NV_NVDLA_CSC_dl_for_check.scala 700:45:@865.4]
  wire [15:0] _T_1850; // @[NV_NVDLA_CSC_dl_for_check.scala 701:42:@868.4]
  wire [15:0] _T_1851; // @[NV_NVDLA_CSC_dl_for_check.scala 701:42:@869.4]
  wire [14:0] _T_1852; // @[NV_NVDLA_CSC_dl_for_check.scala 701:42:@870.4]
  wire  _T_1853; // @[NV_NVDLA_CSC_dl_for_check.scala 702:35:@871.4]
  wire [14:0] _T_1859; // @[NV_NVDLA_CSC_dl_for_check.scala 703:25:@873.4]
  wire [14:0] _T_1860; // @[NV_NVDLA_CSC_dl_for_check.scala 702:25:@874.4]
  wire  _T_1884; // @[Mux.scala 46:19:@884.4]
  wire [12:0] _T_1885; // @[Mux.scala 46:16:@885.4]
  wire  _T_1886; // @[Mux.scala 46:19:@886.4]
  wire [12:0] _T_1887; // @[Mux.scala 46:16:@887.4]
  wire  _T_1888; // @[Mux.scala 46:19:@888.4]
  wire [12:0] _T_1889; // @[Mux.scala 46:16:@889.4]
  wire  _T_1890; // @[Mux.scala 46:19:@890.4]
  wire [12:0] _T_1891; // @[Mux.scala 46:16:@891.4]
  wire [14:0] _GEN_712; // @[NV_NVDLA_CSC_dl_for_check.scala 710:65:@892.4]
  wire  _T_1892; // @[NV_NVDLA_CSC_dl_for_check.scala 710:65:@892.4]
  wire  _T_1893; // @[NV_NVDLA_CSC_dl_for_check.scala 710:85:@893.4]
  wire  _T_1894; // @[NV_NVDLA_CSC_dl_for_check.scala 710:43:@894.4]
  wire  _T_1895; // @[NV_NVDLA_CSC_dl_for_check.scala 712:38:@895.4]
  wire  _T_1897; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@896.4]
  wire  _T_1898; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@897.4]
  wire  _T_1899; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@898.4]
  wire  _T_1902; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@900.4]
  wire  _T_1903; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@901.4]
  wire  _T_1904; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@902.4]
  wire  _T_1907; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@904.4]
  wire  _T_1908; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@905.4]
  wire  _T_1909; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@906.4]
  wire  _T_1912; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@908.4]
  wire  _T_1913; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@909.4]
  wire  _T_1914; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@910.4]
  wire [14:0] _GEN_96; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@916.4]
  wire [14:0] _GEN_97; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@919.4]
  wire [14:0] _GEN_98; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@922.4]
  wire [14:0] _GEN_99; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@925.4]
  wire  _T_1925; // @[NV_NVDLA_CSC_dl_for_check.scala 725:14:@929.4]
  wire [14:0] _GEN_100; // @[NV_NVDLA_CSC_dl_for_check.scala 725:34:@930.4]
  wire [1:0] _GEN_101; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire [1:0] _GEN_102; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire  _GEN_103; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire  _GEN_104; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire  _GEN_106; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire [1:0] _GEN_107; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire  _GEN_108; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire  _GEN_109; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire [8:0] _GEN_110; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  wire [6:0] _T_1935; // @[Cat.scala 30:58:@957.4]
  wire [28:0] _T_1941; // @[Cat.scala 30:58:@963.4]
  reg  _T_1946; // @[NV_NVDLA_CSC_dl_for_check.scala 759:73:@965.4]
  reg [31:0] _RAND_121;
  reg  _T_1949; // @[NV_NVDLA_CSC_dl_for_check.scala 759:73:@966.4]
  reg [31:0] _RAND_122;
  reg  _T_1952; // @[NV_NVDLA_CSC_dl_for_check.scala 759:73:@967.4]
  reg [31:0] _RAND_123;
  reg  _T_1955; // @[NV_NVDLA_CSC_dl_for_check.scala 759:73:@968.4]
  reg [31:0] _RAND_124;
  reg  _T_1958; // @[NV_NVDLA_CSC_dl_for_check.scala 759:73:@969.4]
  reg [31:0] _RAND_125;
  reg  _T_1961; // @[NV_NVDLA_CSC_dl_for_check.scala 759:73:@970.4]
  reg [31:0] _RAND_126;
  reg [28:0] _T_1966; // @[NV_NVDLA_CSC_dl_for_check.scala 761:71:@972.4]
  reg [31:0] _RAND_127;
  reg [28:0] _T_1969; // @[NV_NVDLA_CSC_dl_for_check.scala 761:71:@973.4]
  reg [31:0] _RAND_128;
  reg [28:0] _T_1972; // @[NV_NVDLA_CSC_dl_for_check.scala 761:71:@974.4]
  reg [31:0] _RAND_129;
  reg [28:0] _T_1975; // @[NV_NVDLA_CSC_dl_for_check.scala 761:71:@975.4]
  reg [31:0] _RAND_130;
  reg [28:0] _T_1978; // @[NV_NVDLA_CSC_dl_for_check.scala 761:71:@976.4]
  reg [31:0] _RAND_131;
  reg [28:0] _T_1981; // @[NV_NVDLA_CSC_dl_for_check.scala 761:71:@977.4]
  reg [31:0] _RAND_132;
  wire [28:0] _GEN_111; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1005.4]
  wire [28:0] _GEN_114; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1014.4]
  wire [28:0] _GEN_117; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1023.4]
  wire [28:0] _GEN_120; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1032.4]
  wire [28:0] _GEN_123; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1041.4]
  wire [28:0] _GEN_126; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1050.4]
  wire [1:0] _T_2042; // @[NV_NVDLA_CSC_dl_for_check.scala 794:41:@1058.4]
  wire [1:0] _T_2043; // @[NV_NVDLA_CSC_dl_for_check.scala 795:41:@1059.4]
  wire  _T_2044; // @[NV_NVDLA_CSC_dl_for_check.scala 796:41:@1060.4]
  wire  _T_2045; // @[NV_NVDLA_CSC_dl_for_check.scala 797:42:@1061.4]
  wire [7:0] _T_2046; // @[NV_NVDLA_CSC_dl_for_check.scala 798:41:@1062.4]
  wire [1:0] _T_2047; // @[NV_NVDLA_CSC_dl_for_check.scala 799:45:@1063.4]
  wire  _T_2050; // @[NV_NVDLA_CSC_dl_for_check.scala 802:39:@1066.4]
  wire [8:0] _T_2051; // @[NV_NVDLA_CSC_dl_for_check.scala 803:40:@1067.4]
  reg  _T_2054; // @[NV_NVDLA_CSC_dl_for_check.scala 808:29:@1068.4]
  reg [31:0] _RAND_133;
  reg  _T_2066; // @[NV_NVDLA_CSC_dl_for_check.scala 812:29:@1072.4]
  reg [31:0] _RAND_134;
  reg [511:0] _T_2077; // @[NV_NVDLA_CSC_dl_for_check.scala 817:19:@1076.4]
  reg [511:0] _RAND_135;
  reg [511:0] _T_2085; // @[NV_NVDLA_CSC_dl_for_check.scala 821:19:@1080.4]
  reg [511:0] _RAND_136;
  wire  _T_2108; // @[NV_NVDLA_CSC_dl_for_check.scala 833:69:@1095.4]
  wire  _T_2109; // @[NV_NVDLA_CSC_dl_for_check.scala 833:74:@1096.4]
  wire  _T_2110; // @[NV_NVDLA_CSC_dl_for_check.scala 833:90:@1097.4]
  wire  _T_2111; // @[NV_NVDLA_CSC_dl_for_check.scala 833:88:@1098.4]
  wire  _T_2151; // @[NV_NVDLA_CSC_dl_for_check.scala 848:22:@1132.4]
  wire  _T_2165; // @[NV_NVDLA_CSC_dl_for_check.scala 852:48:@1143.4]
  wire  _T_2166; // @[NV_NVDLA_CSC_dl_for_check.scala 852:22:@1144.4]
  reg [7:0] _T_2185; // @[NV_NVDLA_CSC_dl_for_check.scala 869:29:@1185.4]
  reg [31:0] _RAND_137;
  reg [7:0] _T_2188; // @[NV_NVDLA_CSC_dl_for_check.scala 870:29:@1186.4]
  reg [31:0] _RAND_138;
  reg [7:0] _T_2191; // @[NV_NVDLA_CSC_dl_for_check.scala 871:29:@1187.4]
  reg [31:0] _RAND_139;
  reg [7:0] _T_2194; // @[NV_NVDLA_CSC_dl_for_check.scala 872:29:@1188.4]
  reg [31:0] _RAND_140;
  reg [7:0] _T_2197; // @[NV_NVDLA_CSC_dl_for_check.scala 873:33:@1189.4]
  reg [31:0] _RAND_141;
  reg [7:0] _T_2200; // @[NV_NVDLA_CSC_dl_for_check.scala 874:33:@1190.4]
  reg [31:0] _RAND_142;
  reg [7:0] _T_2203; // @[NV_NVDLA_CSC_dl_for_check.scala 875:33:@1191.4]
  reg [31:0] _RAND_143;
  reg [7:0] _T_2206; // @[NV_NVDLA_CSC_dl_for_check.scala 876:33:@1192.4]
  reg [31:0] _RAND_144;
  reg  _T_2217; // @[NV_NVDLA_CSC_dl_for_check.scala 881:41:@1196.4]
  reg [31:0] _RAND_145;
  reg [26:0] _T_2231; // @[NV_NVDLA_CSC_dl_for_check.scala 883:41:@1201.4]
  reg [31:0] _RAND_146;
  wire [26:0] _T_2243; // @[Cat.scala 30:58:@1211.4]
  wire [26:0] _GEN_137; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1214.4]
  wire [26:0] _GEN_138; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1218.4]
  wire [26:0] _GEN_139; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1222.4]
  wire [26:0] _GEN_140; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1226.4]
  wire  _T_2272; // @[NV_NVDLA_CSC_dl_for_check.scala 909:39:@1252.4]
  wire  _T_2273; // @[NV_NVDLA_CSC_dl_for_check.scala 910:39:@1253.4]
  wire  _T_2274; // @[NV_NVDLA_CSC_dl_for_check.scala 911:39:@1254.4]
  wire  _T_2275; // @[NV_NVDLA_CSC_dl_for_check.scala 912:39:@1255.4]
  wire [8:0] _T_2276; // @[NV_NVDLA_CSC_dl_for_check.scala 914:38:@1256.4]
  wire [8:0] _T_2277; // @[NV_NVDLA_CSC_dl_for_check.scala 915:38:@1257.4]
  wire [8:0] _T_2278; // @[NV_NVDLA_CSC_dl_for_check.scala 916:38:@1258.4]
  wire [8:0] _T_2279; // @[NV_NVDLA_CSC_dl_for_check.scala 917:38:@1259.4]
  wire  _T_2280; // @[NV_NVDLA_CSC_dl_for_check.scala 919:44:@1260.4]
  wire  _T_2281; // @[NV_NVDLA_CSC_dl_for_check.scala 920:44:@1261.4]
  wire  _T_2282; // @[NV_NVDLA_CSC_dl_for_check.scala 921:44:@1262.4]
  wire  _T_2283; // @[NV_NVDLA_CSC_dl_for_check.scala 922:44:@1263.4]
  wire [1:0] _T_2284; // @[NV_NVDLA_CSC_dl_for_check.scala 925:31:@1264.4]
  wire [7:0] _T_2288; // @[NV_NVDLA_CSC_dl_for_check.scala 929:31:@1268.4]
  wire [1:0] _T_2289; // @[NV_NVDLA_CSC_dl_for_check.scala 930:35:@1269.4]
  wire [7:0] _T_2299; // @[NV_NVDLA_CSC_dl_for_check.scala 941:29:@1278.4]
  wire  _T_2310; // @[NV_NVDLA_CSC_dl_for_check.scala 946:50:@1282.4]
  wire [7:0] _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 946:111:@1283.4]
  wire [8:0] _T_2312; // @[NV_NVDLA_CSC_dl_for_check.scala 946:111:@1283.4]
  wire [7:0] _T_2313; // @[NV_NVDLA_CSC_dl_for_check.scala 946:111:@1284.4]
  wire [8:0] _T_2314; // @[NV_NVDLA_CSC_dl_for_check.scala 946:133:@1285.4]
  wire [8:0] _T_2315; // @[NV_NVDLA_CSC_dl_for_check.scala 946:133:@1286.4]
  wire [7:0] _T_2316; // @[NV_NVDLA_CSC_dl_for_check.scala 946:133:@1287.4]
  wire [7:0] _T_2317; // @[NV_NVDLA_CSC_dl_for_check.scala 946:29:@1288.4]
  wire [8:0] _T_2321; // @[NV_NVDLA_CSC_dl_for_check.scala 947:111:@1290.4]
  wire [7:0] _T_2322; // @[NV_NVDLA_CSC_dl_for_check.scala 947:111:@1291.4]
  wire [8:0] _T_2323; // @[NV_NVDLA_CSC_dl_for_check.scala 947:133:@1292.4]
  wire [8:0] _T_2324; // @[NV_NVDLA_CSC_dl_for_check.scala 947:133:@1293.4]
  wire [7:0] _T_2325; // @[NV_NVDLA_CSC_dl_for_check.scala 947:133:@1294.4]
  wire [7:0] _T_2326; // @[NV_NVDLA_CSC_dl_for_check.scala 947:29:@1295.4]
  wire [8:0] _T_2330; // @[NV_NVDLA_CSC_dl_for_check.scala 948:111:@1297.4]
  wire [7:0] _T_2331; // @[NV_NVDLA_CSC_dl_for_check.scala 948:111:@1298.4]
  wire [8:0] _T_2332; // @[NV_NVDLA_CSC_dl_for_check.scala 948:133:@1299.4]
  wire [8:0] _T_2333; // @[NV_NVDLA_CSC_dl_for_check.scala 948:133:@1300.4]
  wire [7:0] _T_2334; // @[NV_NVDLA_CSC_dl_for_check.scala 948:133:@1301.4]
  wire [7:0] _T_2335; // @[NV_NVDLA_CSC_dl_for_check.scala 948:29:@1302.4]
  wire [8:0] _T_2339; // @[NV_NVDLA_CSC_dl_for_check.scala 949:111:@1304.4]
  wire [7:0] _T_2340; // @[NV_NVDLA_CSC_dl_for_check.scala 949:111:@1305.4]
  wire [8:0] _T_2341; // @[NV_NVDLA_CSC_dl_for_check.scala 949:133:@1306.4]
  wire [8:0] _T_2342; // @[NV_NVDLA_CSC_dl_for_check.scala 949:133:@1307.4]
  wire [7:0] _T_2343; // @[NV_NVDLA_CSC_dl_for_check.scala 949:133:@1308.4]
  wire [7:0] _T_2344; // @[NV_NVDLA_CSC_dl_for_check.scala 949:29:@1309.4]
  wire  _T_2346; // @[NV_NVDLA_CSC_dl_for_check.scala 958:52:@1310.4]
  wire  _T_2347; // @[NV_NVDLA_CSC_dl_for_check.scala 958:50:@1311.4]
  wire  _T_2348; // @[NV_NVDLA_CSC_dl_for_check.scala 959:50:@1312.4]
  wire [7:0] _T_2353; // @[NV_NVDLA_CSC_dl_for_check.scala 959:27:@1315.4]
  wire [7:0] _T_2354; // @[NV_NVDLA_CSC_dl_for_check.scala 958:27:@1316.4]
  wire [7:0] _T_2355; // @[NV_NVDLA_CSC_dl_for_check.scala 957:27:@1317.4]
  wire  _T_2357; // @[NV_NVDLA_CSC_dl_for_check.scala 963:52:@1318.4]
  wire  _T_2358; // @[NV_NVDLA_CSC_dl_for_check.scala 963:50:@1319.4]
  wire  _T_2359; // @[NV_NVDLA_CSC_dl_for_check.scala 964:50:@1320.4]
  wire [7:0] _T_2364; // @[NV_NVDLA_CSC_dl_for_check.scala 964:27:@1323.4]
  wire [7:0] _T_2365; // @[NV_NVDLA_CSC_dl_for_check.scala 963:27:@1324.4]
  wire [7:0] _T_2366; // @[NV_NVDLA_CSC_dl_for_check.scala 962:27:@1325.4]
  wire  _T_2368; // @[NV_NVDLA_CSC_dl_for_check.scala 968:52:@1326.4]
  wire  _T_2369; // @[NV_NVDLA_CSC_dl_for_check.scala 968:50:@1327.4]
  wire  _T_2370; // @[NV_NVDLA_CSC_dl_for_check.scala 969:50:@1328.4]
  wire [7:0] _T_2375; // @[NV_NVDLA_CSC_dl_for_check.scala 969:27:@1331.4]
  wire [7:0] _T_2376; // @[NV_NVDLA_CSC_dl_for_check.scala 968:27:@1332.4]
  wire [7:0] _T_2377; // @[NV_NVDLA_CSC_dl_for_check.scala 967:27:@1333.4]
  wire  _T_2379; // @[NV_NVDLA_CSC_dl_for_check.scala 973:52:@1334.4]
  wire  _T_2380; // @[NV_NVDLA_CSC_dl_for_check.scala 973:50:@1335.4]
  wire  _T_2381; // @[NV_NVDLA_CSC_dl_for_check.scala 974:50:@1336.4]
  wire [7:0] _T_2386; // @[NV_NVDLA_CSC_dl_for_check.scala 974:27:@1339.4]
  wire [7:0] _T_2387; // @[NV_NVDLA_CSC_dl_for_check.scala 973:27:@1340.4]
  wire [7:0] _T_2388; // @[NV_NVDLA_CSC_dl_for_check.scala 972:27:@1341.4]
  wire  _T_2389; // @[NV_NVDLA_CSC_dl_for_check.scala 978:46:@1342.4]
  wire  _T_2390; // @[NV_NVDLA_CSC_dl_for_check.scala 978:51:@1343.4]
  wire  _T_2391; // @[NV_NVDLA_CSC_dl_for_check.scala 978:34:@1344.4]
  wire  _T_2392; // @[NV_NVDLA_CSC_dl_for_check.scala 979:46:@1345.4]
  wire  _T_2393; // @[NV_NVDLA_CSC_dl_for_check.scala 979:51:@1346.4]
  wire  _T_2395; // @[NV_NVDLA_CSC_dl_for_check.scala 979:87:@1347.4]
  wire  _T_2396; // @[NV_NVDLA_CSC_dl_for_check.scala 979:69:@1348.4]
  wire  _T_2397; // @[NV_NVDLA_CSC_dl_for_check.scala 979:34:@1349.4]
  wire  _T_2398; // @[NV_NVDLA_CSC_dl_for_check.scala 980:46:@1350.4]
  wire  _T_2399; // @[NV_NVDLA_CSC_dl_for_check.scala 980:51:@1351.4]
  wire  _T_2401; // @[NV_NVDLA_CSC_dl_for_check.scala 980:87:@1352.4]
  wire  _T_2402; // @[NV_NVDLA_CSC_dl_for_check.scala 980:69:@1353.4]
  wire  _T_2403; // @[NV_NVDLA_CSC_dl_for_check.scala 980:34:@1354.4]
  wire  _T_2404; // @[NV_NVDLA_CSC_dl_for_check.scala 981:46:@1355.4]
  wire  _T_2405; // @[NV_NVDLA_CSC_dl_for_check.scala 981:51:@1356.4]
  wire  _T_2408; // @[NV_NVDLA_CSC_dl_for_check.scala 981:69:@1358.4]
  wire  _T_2409; // @[NV_NVDLA_CSC_dl_for_check.scala 981:34:@1359.4]
  wire  _T_2410; // @[NV_NVDLA_CSC_dl_for_check.scala 983:50:@1360.4]
  wire  _T_2411; // @[NV_NVDLA_CSC_dl_for_check.scala 983:55:@1361.4]
  wire  _T_2412; // @[NV_NVDLA_CSC_dl_for_check.scala 983:73:@1362.4]
  wire  _T_2413; // @[NV_NVDLA_CSC_dl_for_check.scala 983:97:@1363.4]
  wire  _T_2414; // @[NV_NVDLA_CSC_dl_for_check.scala 983:38:@1364.4]
  wire  _T_2415; // @[NV_NVDLA_CSC_dl_for_check.scala 984:50:@1365.4]
  wire  _T_2416; // @[NV_NVDLA_CSC_dl_for_check.scala 984:55:@1366.4]
  wire  _T_2417; // @[NV_NVDLA_CSC_dl_for_check.scala 984:73:@1367.4]
  wire  _T_2418; // @[NV_NVDLA_CSC_dl_for_check.scala 984:97:@1368.4]
  wire  _T_2420; // @[NV_NVDLA_CSC_dl_for_check.scala 984:138:@1369.4]
  wire  _T_2421; // @[NV_NVDLA_CSC_dl_for_check.scala 984:120:@1370.4]
  wire  _T_2422; // @[NV_NVDLA_CSC_dl_for_check.scala 984:38:@1371.4]
  wire  _T_2423; // @[NV_NVDLA_CSC_dl_for_check.scala 985:50:@1372.4]
  wire  _T_2424; // @[NV_NVDLA_CSC_dl_for_check.scala 985:55:@1373.4]
  wire  _T_2425; // @[NV_NVDLA_CSC_dl_for_check.scala 985:73:@1374.4]
  wire  _T_2426; // @[NV_NVDLA_CSC_dl_for_check.scala 985:97:@1375.4]
  wire  _T_2428; // @[NV_NVDLA_CSC_dl_for_check.scala 985:138:@1376.4]
  wire  _T_2429; // @[NV_NVDLA_CSC_dl_for_check.scala 985:120:@1377.4]
  wire  _T_2430; // @[NV_NVDLA_CSC_dl_for_check.scala 985:38:@1378.4]
  wire  _T_2431; // @[NV_NVDLA_CSC_dl_for_check.scala 986:50:@1379.4]
  wire  _T_2432; // @[NV_NVDLA_CSC_dl_for_check.scala 986:55:@1380.4]
  wire  _T_2433; // @[NV_NVDLA_CSC_dl_for_check.scala 986:73:@1381.4]
  wire  _T_2434; // @[NV_NVDLA_CSC_dl_for_check.scala 986:97:@1382.4]
  wire  _T_2437; // @[NV_NVDLA_CSC_dl_for_check.scala 986:120:@1384.4]
  wire  _T_2438; // @[NV_NVDLA_CSC_dl_for_check.scala 986:38:@1385.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_dl_for_check.scala 988:24:@1386.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_dl_for_check.scala 989:24:@1389.4]
  wire [7:0] _GEN_143; // @[NV_NVDLA_CSC_dl_for_check.scala 990:24:@1392.4]
  wire [7:0] _GEN_144; // @[NV_NVDLA_CSC_dl_for_check.scala 991:24:@1395.4]
  wire [7:0] _GEN_145; // @[NV_NVDLA_CSC_dl_for_check.scala 992:28:@1398.4]
  wire [7:0] _GEN_146; // @[NV_NVDLA_CSC_dl_for_check.scala 993:28:@1401.4]
  wire [7:0] _GEN_147; // @[NV_NVDLA_CSC_dl_for_check.scala 994:28:@1404.4]
  wire [7:0] _GEN_148; // @[NV_NVDLA_CSC_dl_for_check.scala 995:28:@1407.4]
  wire [7:0] _T_2439; // @[NV_NVDLA_CSC_dl_for_check.scala 1004:55:@1410.4]
  wire [63:0] _T_2442; // @[Cat.scala 30:58:@1413.4]
  wire [127:0] _T_2443; // @[Cat.scala 30:58:@1414.4]
  wire [255:0] _T_2444; // @[Cat.scala 30:58:@1415.4]
  wire [511:0] _T_2445; // @[Cat.scala 30:58:@1416.4]
  wire [511:0] _T_2446; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:23:@1417.4]
  wire [511:0] _T_2450; // @[NV_NVDLA_CSC_dl_for_check.scala 1011:23:@1421.4]
  wire  _T_2456; // @[NV_NVDLA_CSC_dl_for_check.scala 1024:37:@1426.4]
  wire  _T_2459; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:43:@1427.4]
  wire  _T_2460; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:87:@1428.4]
  wire  _T_2462; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:91:@1429.4]
  wire  _T_2463; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:72:@1430.4]
  wire [255:0] _T_2465; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:171:@1431.4]
  wire [511:0] _T_2466; // @[Cat.scala 30:58:@1432.4]
  wire  _T_2472; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:72:@1436.4]
  wire [255:0] _T_2474; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:171:@1437.4]
  wire [511:0] _T_2475; // @[Cat.scala 30:58:@1438.4]
  wire [511:0] _T_2476; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:27:@1439.4]
  wire [511:0] _T_2477; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:27:@1440.4]
  wire [511:0] _T_2478; // @[NV_NVDLA_CSC_dl_for_check.scala 1024:27:@1441.4]
  wire [7:0] _T_2549; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1444.4]
  wire [7:0] _T_2550; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1446.4]
  wire [7:0] _T_2551; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1448.4]
  wire [7:0] _T_2552; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1450.4]
  wire [7:0] _T_2553; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1452.4]
  wire [7:0] _T_2554; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1454.4]
  wire [7:0] _T_2555; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1456.4]
  wire [7:0] _T_2556; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1458.4]
  wire [7:0] _T_2557; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1460.4]
  wire [7:0] _T_2558; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1462.4]
  wire [7:0] _T_2559; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1464.4]
  wire [7:0] _T_2560; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1466.4]
  wire [7:0] _T_2561; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1468.4]
  wire [7:0] _T_2562; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1470.4]
  wire [7:0] _T_2563; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1472.4]
  wire [7:0] _T_2564; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1474.4]
  wire [7:0] _T_2565; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1476.4]
  wire [7:0] _T_2566; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1478.4]
  wire [7:0] _T_2567; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1480.4]
  wire [7:0] _T_2568; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1482.4]
  wire [7:0] _T_2569; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1484.4]
  wire [7:0] _T_2570; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1486.4]
  wire [7:0] _T_2571; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1488.4]
  wire [7:0] _T_2572; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1490.4]
  wire [7:0] _T_2573; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1492.4]
  wire [7:0] _T_2574; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1494.4]
  wire [7:0] _T_2575; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1496.4]
  wire [7:0] _T_2576; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1498.4]
  wire [7:0] _T_2577; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1500.4]
  wire [7:0] _T_2578; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1502.4]
  wire [7:0] _T_2579; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1504.4]
  wire [7:0] _T_2580; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1506.4]
  wire [7:0] _T_2581; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1508.4]
  wire [7:0] _T_2582; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1510.4]
  wire [7:0] _T_2583; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1512.4]
  wire [7:0] _T_2584; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1514.4]
  wire [7:0] _T_2585; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1516.4]
  wire [7:0] _T_2586; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1518.4]
  wire [7:0] _T_2587; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1520.4]
  wire [7:0] _T_2588; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1522.4]
  wire [7:0] _T_2589; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1524.4]
  wire [7:0] _T_2590; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1526.4]
  wire [7:0] _T_2591; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1528.4]
  wire [7:0] _T_2592; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1530.4]
  wire [7:0] _T_2593; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1532.4]
  wire [7:0] _T_2594; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1534.4]
  wire [7:0] _T_2595; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1536.4]
  wire [7:0] _T_2596; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1538.4]
  wire [7:0] _T_2597; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1540.4]
  wire [7:0] _T_2598; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1542.4]
  wire [7:0] _T_2599; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1544.4]
  wire [7:0] _T_2600; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1546.4]
  wire [7:0] _T_2601; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1548.4]
  wire [7:0] _T_2602; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1550.4]
  wire [7:0] _T_2603; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1552.4]
  wire [7:0] _T_2604; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1554.4]
  wire [7:0] _T_2605; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1556.4]
  wire [7:0] _T_2606; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1558.4]
  wire [7:0] _T_2607; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1560.4]
  wire [7:0] _T_2608; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1562.4]
  wire [7:0] _T_2609; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1564.4]
  wire [7:0] _T_2610; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1566.4]
  wire [7:0] _T_2611; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1568.4]
  wire [7:0] _T_2612; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1570.4]
  reg [255:0] _T_2614; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:28:@1572.4]
  reg [255:0] _RAND_147;
  reg [127:0] _T_2616; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:28:@1573.4]
  reg [127:0] _RAND_148;
  reg [127:0] _T_2618; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:28:@1574.4]
  reg [127:0] _RAND_149;
  reg [127:0] _T_2620; // @[NV_NVDLA_CSC_dl_for_check.scala 1050:28:@1575.4]
  reg [127:0] _RAND_150;
  reg [127:0] _T_2622; // @[NV_NVDLA_CSC_dl_for_check.scala 1051:28:@1576.4]
  reg [127:0] _RAND_151;
  reg [127:0] _T_2624; // @[NV_NVDLA_CSC_dl_for_check.scala 1053:28:@1577.4]
  reg [127:0] _RAND_152;
  wire  _T_2625; // @[NV_NVDLA_CSC_dl_for_check.scala 1055:39:@1578.4]
  wire  _T_2626; // @[NV_NVDLA_CSC_dl_for_check.scala 1055:29:@1579.4]
  wire [1023:0] _T_2628; // @[Cat.scala 30:58:@1580.4]
  wire [1023:0] _T_2629; // @[NV_NVDLA_CSC_dl_for_check.scala 1055:28:@1581.4]
  wire  _T_2630; // @[NV_NVDLA_CSC_dl_for_check.scala 1056:39:@1582.4]
  wire  _T_2631; // @[NV_NVDLA_CSC_dl_for_check.scala 1056:29:@1583.4]
  wire [1023:0] _T_2633; // @[Cat.scala 30:58:@1584.4]
  wire [1023:0] _T_2634; // @[NV_NVDLA_CSC_dl_for_check.scala 1056:28:@1585.4]
  wire  _T_2635; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1586.4]
  wire  _T_2636; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:29:@1587.4]
  wire [1023:0] _T_2639; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:28:@1589.4]
  wire  _T_2640; // @[NV_NVDLA_CSC_dl_for_check.scala 1058:39:@1590.4]
  wire  _T_2641; // @[NV_NVDLA_CSC_dl_for_check.scala 1058:29:@1591.4]
  wire [1023:0] _T_2644; // @[NV_NVDLA_CSC_dl_for_check.scala 1058:28:@1593.4]
  wire [10:0] _T_2646; // @[Cat.scala 30:58:@1594.4]
  wire [1023:0] _T_2647; // @[NV_NVDLA_CSC_dl_for_check.scala 1060:41:@1595.4]
  wire [511:0] _T_2648; // @[NV_NVDLA_CSC_dl_for_check.scala 1060:82:@1596.4]
  wire [10:0] _T_2650; // @[Cat.scala 30:58:@1597.4]
  wire [1023:0] _T_2651; // @[NV_NVDLA_CSC_dl_for_check.scala 1061:41:@1598.4]
  wire [511:0] _T_2652; // @[NV_NVDLA_CSC_dl_for_check.scala 1061:82:@1599.4]
  wire [10:0] _T_2654; // @[Cat.scala 30:58:@1600.4]
  wire [1023:0] _T_2655; // @[NV_NVDLA_CSC_dl_for_check.scala 1062:41:@1601.4]
  wire [511:0] _T_2656; // @[NV_NVDLA_CSC_dl_for_check.scala 1062:82:@1602.4]
  wire [10:0] _T_2658; // @[Cat.scala 30:58:@1603.4]
  wire [1023:0] _T_2659; // @[NV_NVDLA_CSC_dl_for_check.scala 1063:41:@1604.4]
  wire [511:0] _T_2660; // @[NV_NVDLA_CSC_dl_for_check.scala 1063:82:@1605.4]
  wire  _T_2661; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:36:@1606.4]
  wire  _T_2662; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:26:@1607.4]
  wire  _T_2665; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:41:@1608.4]
  wire [127:0] _T_2666; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:81:@1609.4]
  wire [511:0] _T_2672; // @[Cat.scala 30:58:@1615.4]
  wire  _T_2674; // @[NV_NVDLA_CSC_dl_for_check.scala 1067:41:@1616.4]
  wire [255:0] _T_2675; // @[NV_NVDLA_CSC_dl_for_check.scala 1067:81:@1617.4]
  wire [511:0] _T_2677; // @[Cat.scala 30:58:@1619.4]
  wire [511:0] _T_2679; // @[NV_NVDLA_CSC_dl_for_check.scala 1067:25:@1621.4]
  wire [511:0] _T_2680; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:25:@1622.4]
  wire [511:0] _T_2681; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:25:@1623.4]
  wire [7:0] _T_2752; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1625.4]
  wire [7:0] _T_2753; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1627.4]
  wire [7:0] _T_2754; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1629.4]
  wire [7:0] _T_2755; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1631.4]
  wire [7:0] _T_2756; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1633.4]
  wire [7:0] _T_2757; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1635.4]
  wire [7:0] _T_2758; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1637.4]
  wire [7:0] _T_2759; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1639.4]
  wire [7:0] _T_2760; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1641.4]
  wire [7:0] _T_2761; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1643.4]
  wire [7:0] _T_2762; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1645.4]
  wire [7:0] _T_2763; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1647.4]
  wire [7:0] _T_2764; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1649.4]
  wire [7:0] _T_2765; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1651.4]
  wire [7:0] _T_2766; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1653.4]
  wire [7:0] _T_2767; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1655.4]
  wire [7:0] _T_2768; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1657.4]
  wire [7:0] _T_2769; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1659.4]
  wire [7:0] _T_2770; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1661.4]
  wire [7:0] _T_2771; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1663.4]
  wire [7:0] _T_2772; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1665.4]
  wire [7:0] _T_2773; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1667.4]
  wire [7:0] _T_2774; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1669.4]
  wire [7:0] _T_2775; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1671.4]
  wire [7:0] _T_2776; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1673.4]
  wire [7:0] _T_2777; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1675.4]
  wire [7:0] _T_2778; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1677.4]
  wire [7:0] _T_2779; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1679.4]
  wire [7:0] _T_2780; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1681.4]
  wire [7:0] _T_2781; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1683.4]
  wire [7:0] _T_2782; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1685.4]
  wire [7:0] _T_2783; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1687.4]
  wire [7:0] _T_2784; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1689.4]
  wire [7:0] _T_2785; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1691.4]
  wire [7:0] _T_2786; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1693.4]
  wire [7:0] _T_2787; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1695.4]
  wire [7:0] _T_2788; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1697.4]
  wire [7:0] _T_2789; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1699.4]
  wire [7:0] _T_2790; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1701.4]
  wire [7:0] _T_2791; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1703.4]
  wire [7:0] _T_2792; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1705.4]
  wire [7:0] _T_2793; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1707.4]
  wire [7:0] _T_2794; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1709.4]
  wire [7:0] _T_2795; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1711.4]
  wire [7:0] _T_2796; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1713.4]
  wire [7:0] _T_2797; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1715.4]
  wire [7:0] _T_2798; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1717.4]
  wire [7:0] _T_2799; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1719.4]
  wire [7:0] _T_2800; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1721.4]
  wire [7:0] _T_2801; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1723.4]
  wire [7:0] _T_2802; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1725.4]
  wire [7:0] _T_2803; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1727.4]
  wire [7:0] _T_2804; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1729.4]
  wire [7:0] _T_2805; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1731.4]
  wire [7:0] _T_2806; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1733.4]
  wire [7:0] _T_2807; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1735.4]
  wire [7:0] _T_2808; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1737.4]
  wire [7:0] _T_2809; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1739.4]
  wire [7:0] _T_2810; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1741.4]
  wire [7:0] _T_2811; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1743.4]
  wire [7:0] _T_2812; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1745.4]
  wire [7:0] _T_2813; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1747.4]
  wire [7:0] _T_2814; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1749.4]
  wire [7:0] _T_2815; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1751.4]
  wire  _T_2817; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:59:@1753.4]
  wire  _T_2818; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:41:@1754.4]
  wire  _T_2820; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:59:@1755.4]
  wire  _T_2821; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:41:@1756.4]
  wire  _T_2824; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:41:@1758.4]
  wire [511:0] _GEN_149; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:24:@1759.4]
  wire [255:0] _GEN_150; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:24:@1762.4]
  wire [511:0] _GEN_151; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:24:@1762.4]
  wire [511:0] _GEN_154; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:24:@1766.4]
  wire [318:0] _T_2830; // @[NV_NVDLA_CSC_dl_for_check.scala 1096:56:@1772.4]
  wire [63:0] _T_2831; // @[NV_NVDLA_CSC_dl_for_check.scala 1096:73:@1773.4]
  wire [63:0] _T_2832; // @[NV_NVDLA_CSC_dl_for_check.scala 1096:24:@1774.4]
  wire  _T_2834; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:51:@1775.4]
  wire [63:0] _T_2841; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:32:@1777.4]
  wire  _T_2843; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:51:@1778.4]
  wire [31:0] _T_2850; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:32:@1780.4]
  wire  _T_2852; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:51:@1781.4]
  wire [31:0] _T_2859; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:32:@1783.4]
  wire [31:0] _T_2860; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:57:@1784.4]
  wire [63:0] _T_2866; // @[Cat.scala 30:58:@1786.4]
  wire [15:0] _T_2867; // @[NV_NVDLA_CSC_dl_for_check.scala 1103:57:@1787.4]
  wire [15:0] _T_2868; // @[NV_NVDLA_CSC_dl_for_check.scala 1103:106:@1788.4]
  wire [15:0] _T_2869; // @[NV_NVDLA_CSC_dl_for_check.scala 1103:155:@1789.4]
  wire [63:0] _T_2877; // @[Cat.scala 30:58:@1793.4]
  wire  _T_2879; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:43:@1794.4]
  wire [15:0] _T_2880; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:89:@1795.4]
  wire [63:0] _T_2882; // @[Cat.scala 30:58:@1797.4]
  wire [63:0] _T_2883; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:116:@1798.4]
  wire  _T_2885; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:43:@1799.4]
  wire [31:0] _T_2886; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:89:@1800.4]
  wire [63:0] _T_2887; // @[Cat.scala 30:58:@1801.4]
  wire [63:0] _T_2888; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:116:@1802.4]
  wire [63:0] _T_2889; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:26:@1803.4]
  wire [63:0] _T_2890; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:26:@1804.4]
  wire  _T_2891; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:35:@1805.4]
  wire [7:0] _T_2892_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire [7:0] _T_2892_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  wire  _T_3025; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1807.4]
  wire  _T_3027; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1808.4]
  wire  _T_3029; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1809.4]
  wire  _T_3031; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1810.4]
  wire  _T_3033; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1811.4]
  wire  _T_3035; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1812.4]
  wire  _T_3037; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1813.4]
  wire  _T_3039; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1814.4]
  wire  _T_3041; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1815.4]
  wire  _T_3043; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1816.4]
  wire  _T_3045; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1817.4]
  wire  _T_3047; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1818.4]
  wire  _T_3049; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1819.4]
  wire  _T_3051; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1820.4]
  wire  _T_3053; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1821.4]
  wire  _T_3055; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1822.4]
  wire  _T_3057; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1823.4]
  wire  _T_3059; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1824.4]
  wire  _T_3061; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1825.4]
  wire  _T_3063; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1826.4]
  wire  _T_3065; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1827.4]
  wire  _T_3067; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1828.4]
  wire  _T_3069; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1829.4]
  wire  _T_3071; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1830.4]
  wire  _T_3073; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1831.4]
  wire  _T_3075; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1832.4]
  wire  _T_3077; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1833.4]
  wire  _T_3079; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1834.4]
  wire  _T_3081; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1835.4]
  wire  _T_3083; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1836.4]
  wire  _T_3085; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1837.4]
  wire  _T_3087; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1838.4]
  wire  _T_3089; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1839.4]
  wire  _T_3091; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1840.4]
  wire  _T_3093; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1841.4]
  wire  _T_3095; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1842.4]
  wire  _T_3097; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1843.4]
  wire  _T_3099; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1844.4]
  wire  _T_3101; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1845.4]
  wire  _T_3103; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1846.4]
  wire  _T_3105; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1847.4]
  wire  _T_3107; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1848.4]
  wire  _T_3109; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1849.4]
  wire  _T_3111; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1850.4]
  wire  _T_3113; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1851.4]
  wire  _T_3115; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1852.4]
  wire  _T_3117; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1853.4]
  wire  _T_3119; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1854.4]
  wire  _T_3121; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1855.4]
  wire  _T_3123; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1856.4]
  wire  _T_3125; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1857.4]
  wire  _T_3127; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1858.4]
  wire  _T_3129; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1859.4]
  wire  _T_3131; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1860.4]
  wire  _T_3133; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1861.4]
  wire  _T_3135; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1862.4]
  wire  _T_3137; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1863.4]
  wire  _T_3139; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1864.4]
  wire  _T_3141; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1865.4]
  wire  _T_3143; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1866.4]
  wire  _T_3145; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1867.4]
  wire  _T_3147; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1868.4]
  wire  _T_3149; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1869.4]
  wire  _T_3151; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1870.4]
  wire  _T_3222; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1936.4]
  wire  _T_3223; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1937.4]
  wire  _T_3224; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1938.4]
  wire  _T_3225; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1939.4]
  wire  _T_3226; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1940.4]
  wire  _T_3227; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1941.4]
  wire  _T_3228; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1942.4]
  wire  _T_3229; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1943.4]
  wire  _T_3230; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1944.4]
  wire  _T_3231; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1945.4]
  wire  _T_3232; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1946.4]
  wire  _T_3233; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1947.4]
  wire  _T_3234; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1948.4]
  wire  _T_3235; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1949.4]
  wire  _T_3236; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1950.4]
  wire  _T_3237; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1951.4]
  wire  _T_3238; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1952.4]
  wire  _T_3239; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1953.4]
  wire  _T_3240; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1954.4]
  wire  _T_3241; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1955.4]
  wire  _T_3242; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1956.4]
  wire  _T_3243; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1957.4]
  wire  _T_3244; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1958.4]
  wire  _T_3245; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1959.4]
  wire  _T_3246; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1960.4]
  wire  _T_3247; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1961.4]
  wire  _T_3248; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1962.4]
  wire  _T_3249; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1963.4]
  wire  _T_3250; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1964.4]
  wire  _T_3251; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1965.4]
  wire  _T_3252; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1966.4]
  wire  _T_3253; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1967.4]
  wire  _T_3254; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1968.4]
  wire  _T_3255; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1969.4]
  wire  _T_3256; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1970.4]
  wire  _T_3257; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1971.4]
  wire  _T_3258; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1972.4]
  wire  _T_3259; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1973.4]
  wire  _T_3260; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1974.4]
  wire  _T_3261; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1975.4]
  wire  _T_3262; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1976.4]
  wire  _T_3263; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1977.4]
  wire  _T_3264; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1978.4]
  wire  _T_3265; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1979.4]
  wire  _T_3266; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1980.4]
  wire  _T_3267; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1981.4]
  wire  _T_3268; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1982.4]
  wire  _T_3269; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1983.4]
  wire  _T_3270; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1984.4]
  wire  _T_3271; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1985.4]
  wire  _T_3272; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1986.4]
  wire  _T_3273; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1987.4]
  wire  _T_3274; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1988.4]
  wire  _T_3275; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1989.4]
  wire  _T_3276; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1990.4]
  wire  _T_3277; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1991.4]
  wire  _T_3278; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1992.4]
  wire  _T_3279; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1993.4]
  wire  _T_3280; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1994.4]
  wire  _T_3281; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1995.4]
  wire  _T_3282; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1996.4]
  wire  _T_3283; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1997.4]
  wire  _T_3284; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1998.4]
  wire  _T_3285; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1999.4]
  wire  _T_3286; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2000.4]
  wire  _T_3287; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2001.4]
  wire  _T_3288; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2002.4]
  wire  _T_3289; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2003.4]
  wire  _T_3290; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2004.4]
  wire  _T_3291; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2005.4]
  wire  _T_3292; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2006.4]
  wire  _T_3293; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2007.4]
  wire  _T_3294; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2008.4]
  wire  _T_3295; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2009.4]
  wire  _T_3296; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2010.4]
  wire  _T_3297; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2011.4]
  wire  _T_3298; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2012.4]
  wire  _T_3299; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2013.4]
  wire  _T_3300; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2014.4]
  wire  _T_3301; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2015.4]
  wire  _T_3302; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2016.4]
  wire  _T_3303; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2017.4]
  wire  _T_3304; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2018.4]
  wire  _T_3305; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2019.4]
  wire  _T_3306; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2020.4]
  wire  _T_3307; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2021.4]
  wire  _T_3308; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2022.4]
  wire  _T_3309; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2023.4]
  wire  _T_3310; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2024.4]
  wire  _T_3311; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2025.4]
  wire  _T_3312; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2026.4]
  wire  _T_3313; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2027.4]
  wire  _T_3314; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2028.4]
  wire  _T_3315; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2029.4]
  wire  _T_3316; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2030.4]
  wire  _T_3317; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2031.4]
  wire  _T_3318; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2032.4]
  wire  _T_3319; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2033.4]
  wire  _T_3320; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2034.4]
  wire  _T_3321; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2035.4]
  wire  _T_3322; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2036.4]
  wire  _T_3323; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2037.4]
  wire  _T_3324; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2038.4]
  wire  _T_3325; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2039.4]
  wire  _T_3326; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2040.4]
  wire  _T_3327; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2041.4]
  wire  _T_3328; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2042.4]
  wire  _T_3329; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2043.4]
  wire  _T_3330; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2044.4]
  wire  _T_3331; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2045.4]
  wire  _T_3332; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2046.4]
  wire  _T_3333; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2047.4]
  wire  _T_3334; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2048.4]
  wire  _T_3335; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2049.4]
  wire  _T_3336; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2050.4]
  wire  _T_3337; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2051.4]
  wire  _T_3338; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2052.4]
  wire  _T_3339; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2053.4]
  wire  _T_3340; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2054.4]
  wire  _T_3341; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2055.4]
  wire  _T_3342; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2056.4]
  wire  _T_3343; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2057.4]
  wire  _T_3344; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2058.4]
  wire  _T_3345; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2059.4]
  wire  _T_3346; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2060.4]
  wire  _T_3347; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2061.4]
  wire  _T_3348; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2062.4]
  wire  _T_3349; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2063.4]
  reg  _T_3422; // @[NV_NVDLA_CSC_dl_for_check.scala 1119:27:@2129.4]
  reg [31:0] _RAND_153;
  reg  _T_3692_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_154;
  reg  _T_3692_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_155;
  reg  _T_3692_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_156;
  reg  _T_3692_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_157;
  reg  _T_3692_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_158;
  reg  _T_3692_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_159;
  reg  _T_3692_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_160;
  reg  _T_3692_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_161;
  reg  _T_3692_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_162;
  reg  _T_3692_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_163;
  reg  _T_3692_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_164;
  reg  _T_3692_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_165;
  reg  _T_3692_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_166;
  reg  _T_3692_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_167;
  reg  _T_3692_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_168;
  reg  _T_3692_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_169;
  reg  _T_3692_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_170;
  reg  _T_3692_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_171;
  reg  _T_3692_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_172;
  reg  _T_3692_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_173;
  reg  _T_3692_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_174;
  reg  _T_3692_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_175;
  reg  _T_3692_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_176;
  reg  _T_3692_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_177;
  reg  _T_3692_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_178;
  reg  _T_3692_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_179;
  reg  _T_3692_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_180;
  reg  _T_3692_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_181;
  reg  _T_3692_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_182;
  reg  _T_3692_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_183;
  reg  _T_3692_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_184;
  reg  _T_3692_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_185;
  reg  _T_3692_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_186;
  reg  _T_3692_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_187;
  reg  _T_3692_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_188;
  reg  _T_3692_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_189;
  reg  _T_3692_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_190;
  reg  _T_3692_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_191;
  reg  _T_3692_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_192;
  reg  _T_3692_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_193;
  reg  _T_3692_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_194;
  reg  _T_3692_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_195;
  reg  _T_3692_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_196;
  reg  _T_3692_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_197;
  reg  _T_3692_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_198;
  reg  _T_3692_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_199;
  reg  _T_3692_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_200;
  reg  _T_3692_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_201;
  reg  _T_3692_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_202;
  reg  _T_3692_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_203;
  reg  _T_3692_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_204;
  reg  _T_3692_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_205;
  reg  _T_3692_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_206;
  reg  _T_3692_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_207;
  reg  _T_3692_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_208;
  reg  _T_3692_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_209;
  reg  _T_3692_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_210;
  reg  _T_3692_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_211;
  reg  _T_3692_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_212;
  reg  _T_3692_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_213;
  reg  _T_3692_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_214;
  reg  _T_3692_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_215;
  reg  _T_3692_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_216;
  reg  _T_3692_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:34:@2196.4]
  reg [31:0] _RAND_217;
  reg [7:0] _T_3892_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_218;
  reg [7:0] _T_3892_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_219;
  reg [7:0] _T_3892_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_220;
  reg [7:0] _T_3892_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_221;
  reg [7:0] _T_3892_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_222;
  reg [7:0] _T_3892_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_223;
  reg [7:0] _T_3892_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_224;
  reg [7:0] _T_3892_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_225;
  reg [7:0] _T_3892_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_226;
  reg [7:0] _T_3892_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_227;
  reg [7:0] _T_3892_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_228;
  reg [7:0] _T_3892_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_229;
  reg [7:0] _T_3892_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_230;
  reg [7:0] _T_3892_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_231;
  reg [7:0] _T_3892_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_232;
  reg [7:0] _T_3892_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_233;
  reg [7:0] _T_3892_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_234;
  reg [7:0] _T_3892_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_235;
  reg [7:0] _T_3892_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_236;
  reg [7:0] _T_3892_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_237;
  reg [7:0] _T_3892_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_238;
  reg [7:0] _T_3892_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_239;
  reg [7:0] _T_3892_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_240;
  reg [7:0] _T_3892_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_241;
  reg [7:0] _T_3892_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_242;
  reg [7:0] _T_3892_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_243;
  reg [7:0] _T_3892_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_244;
  reg [7:0] _T_3892_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_245;
  reg [7:0] _T_3892_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_246;
  reg [7:0] _T_3892_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_247;
  reg [7:0] _T_3892_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_248;
  reg [7:0] _T_3892_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_249;
  reg [7:0] _T_3892_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_250;
  reg [7:0] _T_3892_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_251;
  reg [7:0] _T_3892_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_252;
  reg [7:0] _T_3892_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_253;
  reg [7:0] _T_3892_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_254;
  reg [7:0] _T_3892_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_255;
  reg [7:0] _T_3892_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_256;
  reg [7:0] _T_3892_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_257;
  reg [7:0] _T_3892_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_258;
  reg [7:0] _T_3892_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_259;
  reg [7:0] _T_3892_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_260;
  reg [7:0] _T_3892_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_261;
  reg [7:0] _T_3892_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_262;
  reg [7:0] _T_3892_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_263;
  reg [7:0] _T_3892_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_264;
  reg [7:0] _T_3892_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_265;
  reg [7:0] _T_3892_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_266;
  reg [7:0] _T_3892_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_267;
  reg [7:0] _T_3892_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_268;
  reg [7:0] _T_3892_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_269;
  reg [7:0] _T_3892_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_270;
  reg [7:0] _T_3892_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_271;
  reg [7:0] _T_3892_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_272;
  reg [7:0] _T_3892_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_273;
  reg [7:0] _T_3892_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_274;
  reg [7:0] _T_3892_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_275;
  reg [7:0] _T_3892_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_276;
  reg [7:0] _T_3892_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_277;
  reg [7:0] _T_3892_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_278;
  reg [7:0] _T_3892_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_279;
  reg [7:0] _T_3892_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_280;
  reg [7:0] _T_3892_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:30:@2197.4]
  reg [31:0] _RAND_281;
  wire  _GEN_156; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_209; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  wire  _T_3959; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2268.4]
  wire  _T_3960; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2272.4]
  wire  _T_3961; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2276.4]
  wire  _T_3962; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2280.4]
  wire  _T_3963; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2284.4]
  wire  _T_3964; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2288.4]
  wire  _T_3965; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2292.4]
  wire  _T_3966; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2296.4]
  wire  _T_3967; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2300.4]
  wire  _T_3968; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2304.4]
  wire  _T_3969; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2308.4]
  wire  _T_3970; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2312.4]
  wire  _T_3971; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2316.4]
  wire  _T_3972; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2320.4]
  wire  _T_3973; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2324.4]
  wire  _T_3974; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2328.4]
  wire  _T_3975; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2332.4]
  wire  _T_3976; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2336.4]
  wire  _T_3977; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2340.4]
  wire  _T_3978; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2344.4]
  wire  _T_3979; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2348.4]
  wire  _T_3980; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2352.4]
  wire  _T_3981; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2356.4]
  wire  _T_3982; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2360.4]
  wire  _T_3983; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2364.4]
  wire  _T_3984; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2368.4]
  wire  _T_3985; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2372.4]
  wire  _T_3986; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2376.4]
  wire  _T_3987; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2380.4]
  wire  _T_3988; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2384.4]
  wire  _T_3989; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2388.4]
  wire  _T_3990; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2392.4]
  wire  _T_3991; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2396.4]
  wire  _T_3992; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2400.4]
  wire  _T_3993; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2404.4]
  wire  _T_3994; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2408.4]
  wire  _T_3995; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2412.4]
  wire  _T_3996; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2416.4]
  wire  _T_3997; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2420.4]
  wire  _T_3998; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2424.4]
  wire  _T_3999; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2428.4]
  wire  _T_4000; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2432.4]
  wire  _T_4001; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2436.4]
  wire  _T_4002; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2440.4]
  wire  _T_4003; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2444.4]
  wire  _T_4004; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2448.4]
  wire  _T_4005; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2452.4]
  wire  _T_4006; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2456.4]
  wire  _T_4007; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2460.4]
  wire  _T_4008; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2464.4]
  wire  _T_4009; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2468.4]
  wire  _T_4010; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2472.4]
  wire  _T_4011; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2476.4]
  wire  _T_4012; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2480.4]
  wire  _T_4013; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2484.4]
  wire  _T_4014; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2488.4]
  wire  _T_4015; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2492.4]
  wire  _T_4016; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2496.4]
  wire  _T_4017; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2500.4]
  wire  _T_4018; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2504.4]
  wire  _T_4019; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2508.4]
  wire  _T_4020; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2512.4]
  wire  _T_4021; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2516.4]
  wire  _T_4022; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2520.4]
  reg  _T_4025; // @[NV_NVDLA_CSC_dl_for_check.scala 1147:26:@2524.4]
  reg [31:0] _RAND_282;
  reg  _T_4292_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_283;
  reg  _T_4292_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_284;
  reg  _T_4292_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_285;
  reg  _T_4292_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_286;
  reg  _T_4292_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_287;
  reg  _T_4292_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_288;
  reg  _T_4292_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_289;
  reg  _T_4292_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_290;
  reg  _T_4292_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_291;
  reg  _T_4292_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_292;
  reg  _T_4292_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_293;
  reg  _T_4292_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_294;
  reg  _T_4292_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_295;
  reg  _T_4292_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_296;
  reg  _T_4292_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_297;
  reg  _T_4292_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_298;
  reg  _T_4292_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_299;
  reg  _T_4292_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_300;
  reg  _T_4292_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_301;
  reg  _T_4292_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_302;
  reg  _T_4292_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_303;
  reg  _T_4292_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_304;
  reg  _T_4292_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_305;
  reg  _T_4292_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_306;
  reg  _T_4292_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_307;
  reg  _T_4292_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_308;
  reg  _T_4292_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_309;
  reg  _T_4292_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_310;
  reg  _T_4292_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_311;
  reg  _T_4292_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_312;
  reg  _T_4292_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_313;
  reg  _T_4292_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_314;
  reg  _T_4292_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_315;
  reg  _T_4292_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_316;
  reg  _T_4292_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_317;
  reg  _T_4292_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_318;
  reg  _T_4292_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_319;
  reg  _T_4292_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_320;
  reg  _T_4292_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_321;
  reg  _T_4292_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_322;
  reg  _T_4292_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_323;
  reg  _T_4292_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_324;
  reg  _T_4292_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_325;
  reg  _T_4292_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_326;
  reg  _T_4292_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_327;
  reg  _T_4292_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_328;
  reg  _T_4292_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_329;
  reg  _T_4292_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_330;
  reg  _T_4292_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_331;
  reg  _T_4292_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_332;
  reg  _T_4292_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_333;
  reg  _T_4292_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_334;
  reg  _T_4292_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_335;
  reg  _T_4292_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_336;
  reg  _T_4292_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_337;
  reg  _T_4292_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_338;
  reg  _T_4292_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_339;
  reg  _T_4292_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_340;
  reg  _T_4292_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_341;
  reg  _T_4292_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_342;
  reg  _T_4292_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_343;
  reg  _T_4292_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_344;
  reg  _T_4292_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_345;
  reg  _T_4292_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:26:@2590.4]
  reg [31:0] _RAND_346;
  reg [8:0] _T_4491; // @[NV_NVDLA_CSC_dl_for_check.scala 1149:26:@2591.4]
  reg [31:0] _RAND_347;
  reg [7:0] _T_4495_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_348;
  reg [7:0] _T_4495_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_349;
  reg [7:0] _T_4495_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_350;
  reg [7:0] _T_4495_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_351;
  reg [7:0] _T_4495_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_352;
  reg [7:0] _T_4495_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_353;
  reg [7:0] _T_4495_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_354;
  reg [7:0] _T_4495_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_355;
  reg [7:0] _T_4495_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_356;
  reg [7:0] _T_4495_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_357;
  reg [7:0] _T_4495_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_358;
  reg [7:0] _T_4495_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_359;
  reg [7:0] _T_4495_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_360;
  reg [7:0] _T_4495_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_361;
  reg [7:0] _T_4495_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_362;
  reg [7:0] _T_4495_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_363;
  reg [7:0] _T_4495_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_364;
  reg [7:0] _T_4495_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_365;
  reg [7:0] _T_4495_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_366;
  reg [7:0] _T_4495_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_367;
  reg [7:0] _T_4495_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_368;
  reg [7:0] _T_4495_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_369;
  reg [7:0] _T_4495_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_370;
  reg [7:0] _T_4495_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_371;
  reg [7:0] _T_4495_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_372;
  reg [7:0] _T_4495_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_373;
  reg [7:0] _T_4495_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_374;
  reg [7:0] _T_4495_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_375;
  reg [7:0] _T_4495_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_376;
  reg [7:0] _T_4495_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_377;
  reg [7:0] _T_4495_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_378;
  reg [7:0] _T_4495_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_379;
  reg [7:0] _T_4495_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_380;
  reg [7:0] _T_4495_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_381;
  reg [7:0] _T_4495_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_382;
  reg [7:0] _T_4495_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_383;
  reg [7:0] _T_4495_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_384;
  reg [7:0] _T_4495_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_385;
  reg [7:0] _T_4495_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_386;
  reg [7:0] _T_4495_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_387;
  reg [7:0] _T_4495_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_388;
  reg [7:0] _T_4495_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_389;
  reg [7:0] _T_4495_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_390;
  reg [7:0] _T_4495_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_391;
  reg [7:0] _T_4495_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_392;
  reg [7:0] _T_4495_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_393;
  reg [7:0] _T_4495_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_394;
  reg [7:0] _T_4495_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_395;
  reg [7:0] _T_4495_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_396;
  reg [7:0] _T_4495_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_397;
  reg [7:0] _T_4495_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_398;
  reg [7:0] _T_4495_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_399;
  reg [7:0] _T_4495_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_400;
  reg [7:0] _T_4495_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_401;
  reg [7:0] _T_4495_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_402;
  reg [7:0] _T_4495_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_403;
  reg [7:0] _T_4495_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_404;
  reg [7:0] _T_4495_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_405;
  reg [7:0] _T_4495_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_406;
  reg [7:0] _T_4495_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_407;
  reg [7:0] _T_4495_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_408;
  reg [7:0] _T_4495_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_409;
  reg [7:0] _T_4495_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_410;
  reg [7:0] _T_4495_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1150:22:@2592.4]
  reg [31:0] _RAND_411;
  wire  _T_4562; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:24:@2593.4]
  wire  _T_4697_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4697_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  wire  _T_4829; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:19:@2661.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_289; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  wire [8:0] _GEN_348; // @[NV_NVDLA_CSC_dl_for_check.scala 1160:19:@2728.4]
  reg  _T_4832; // @[NV_NVDLA_CSC_dl_for_check.scala 1173:29:@2923.4]
  reg [31:0] _RAND_412;
  wire  _T_4833; // @[NV_NVDLA_CSC_dl_for_check.scala 1174:27:@2925.4]
  wire [8:0] _T_4835; // @[NV_NVDLA_CSC_dl_for_check.scala 1174:26:@2926.4]
  reg  _T_4838; // @[NV_NVDLA_CSC_dl_for_check.scala 1176:33:@2927.4]
  reg [31:0] _RAND_413;
  reg  _T_4841; // @[NV_NVDLA_CSC_dl_for_check.scala 1177:33:@2930.4]
  reg [31:0] _RAND_414;
  wire  _T_4843; // @[NV_NVDLA_CSC_dl_for_check.scala 1178:85:@2933.4]
  reg [8:0] _T_4845; // @[Reg.scala 19:20:@2934.4]
  reg [31:0] _RAND_415;
  wire [8:0] _GEN_413; // @[Reg.scala 20:19:@2935.4]
  reg [8:0] _T_4849; // @[Reg.scala 19:20:@2940.4]
  reg [31:0] _RAND_416;
  wire [8:0] _GEN_414; // @[Reg.scala 20:19:@2941.4]
  reg  _T_5117_0; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_417;
  reg  _T_5117_1; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_418;
  reg  _T_5117_2; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_419;
  reg  _T_5117_3; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_420;
  reg  _T_5117_4; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_421;
  reg  _T_5117_5; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_422;
  reg  _T_5117_6; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_423;
  reg  _T_5117_7; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_424;
  reg  _T_5117_8; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_425;
  reg  _T_5117_9; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_426;
  reg  _T_5117_10; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_427;
  reg  _T_5117_11; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_428;
  reg  _T_5117_12; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_429;
  reg  _T_5117_13; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_430;
  reg  _T_5117_14; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_431;
  reg  _T_5117_15; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_432;
  reg  _T_5117_16; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_433;
  reg  _T_5117_17; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_434;
  reg  _T_5117_18; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_435;
  reg  _T_5117_19; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_436;
  reg  _T_5117_20; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_437;
  reg  _T_5117_21; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_438;
  reg  _T_5117_22; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_439;
  reg  _T_5117_23; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_440;
  reg  _T_5117_24; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_441;
  reg  _T_5117_25; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_442;
  reg  _T_5117_26; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_443;
  reg  _T_5117_27; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_444;
  reg  _T_5117_28; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_445;
  reg  _T_5117_29; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_446;
  reg  _T_5117_30; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_447;
  reg  _T_5117_31; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_448;
  reg  _T_5117_32; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_449;
  reg  _T_5117_33; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_450;
  reg  _T_5117_34; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_451;
  reg  _T_5117_35; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_452;
  reg  _T_5117_36; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_453;
  reg  _T_5117_37; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_454;
  reg  _T_5117_38; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_455;
  reg  _T_5117_39; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_456;
  reg  _T_5117_40; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_457;
  reg  _T_5117_41; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_458;
  reg  _T_5117_42; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_459;
  reg  _T_5117_43; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_460;
  reg  _T_5117_44; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_461;
  reg  _T_5117_45; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_462;
  reg  _T_5117_46; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_463;
  reg  _T_5117_47; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_464;
  reg  _T_5117_48; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_465;
  reg  _T_5117_49; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_466;
  reg  _T_5117_50; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_467;
  reg  _T_5117_51; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_468;
  reg  _T_5117_52; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_469;
  reg  _T_5117_53; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_470;
  reg  _T_5117_54; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_471;
  reg  _T_5117_55; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_472;
  reg  _T_5117_56; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_473;
  reg  _T_5117_57; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_474;
  reg  _T_5117_58; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_475;
  reg  _T_5117_59; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_476;
  reg  _T_5117_60; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_477;
  reg  _T_5117_61; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_478;
  reg  _T_5117_62; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_479;
  reg  _T_5117_63; // @[Reg.scala 19:20:@3011.4]
  reg [31:0] _RAND_480;
  wire  _GEN_415; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_416; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_417; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_418; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_419; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_420; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_421; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_422; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_423; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_424; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_425; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_426; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_427; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_428; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_429; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_430; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_431; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_432; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_433; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_434; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_435; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_436; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_437; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_438; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_439; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_440; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_441; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_442; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_443; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_444; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_445; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_446; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_447; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_448; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_449; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_450; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_451; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_452; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_453; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_454; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_455; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_456; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_457; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_458; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_459; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_460; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_461; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_462; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_463; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_464; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_465; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_466; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_467; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_468; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_469; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_470; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_471; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_472; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_473; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_474; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_475; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_476; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_477; // @[Reg.scala 20:19:@3012.4]
  wire  _GEN_478; // @[Reg.scala 20:19:@3012.4]
  reg  _T_5581_0; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_481;
  reg  _T_5581_1; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_482;
  reg  _T_5581_2; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_483;
  reg  _T_5581_3; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_484;
  reg  _T_5581_4; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_485;
  reg  _T_5581_5; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_486;
  reg  _T_5581_6; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_487;
  reg  _T_5581_7; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_488;
  reg  _T_5581_8; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_489;
  reg  _T_5581_9; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_490;
  reg  _T_5581_10; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_491;
  reg  _T_5581_11; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_492;
  reg  _T_5581_12; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_493;
  reg  _T_5581_13; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_494;
  reg  _T_5581_14; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_495;
  reg  _T_5581_15; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_496;
  reg  _T_5581_16; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_497;
  reg  _T_5581_17; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_498;
  reg  _T_5581_18; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_499;
  reg  _T_5581_19; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_500;
  reg  _T_5581_20; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_501;
  reg  _T_5581_21; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_502;
  reg  _T_5581_22; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_503;
  reg  _T_5581_23; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_504;
  reg  _T_5581_24; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_505;
  reg  _T_5581_25; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_506;
  reg  _T_5581_26; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_507;
  reg  _T_5581_27; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_508;
  reg  _T_5581_28; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_509;
  reg  _T_5581_29; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_510;
  reg  _T_5581_30; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_511;
  reg  _T_5581_31; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_512;
  reg  _T_5581_32; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_513;
  reg  _T_5581_33; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_514;
  reg  _T_5581_34; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_515;
  reg  _T_5581_35; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_516;
  reg  _T_5581_36; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_517;
  reg  _T_5581_37; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_518;
  reg  _T_5581_38; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_519;
  reg  _T_5581_39; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_520;
  reg  _T_5581_40; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_521;
  reg  _T_5581_41; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_522;
  reg  _T_5581_42; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_523;
  reg  _T_5581_43; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_524;
  reg  _T_5581_44; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_525;
  reg  _T_5581_45; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_526;
  reg  _T_5581_46; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_527;
  reg  _T_5581_47; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_528;
  reg  _T_5581_48; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_529;
  reg  _T_5581_49; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_530;
  reg  _T_5581_50; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_531;
  reg  _T_5581_51; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_532;
  reg  _T_5581_52; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_533;
  reg  _T_5581_53; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_534;
  reg  _T_5581_54; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_535;
  reg  _T_5581_55; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_536;
  reg  _T_5581_56; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_537;
  reg  _T_5581_57; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_538;
  reg  _T_5581_58; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_539;
  reg  _T_5581_59; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_540;
  reg  _T_5581_60; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_541;
  reg  _T_5581_61; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_542;
  reg  _T_5581_62; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_543;
  reg  _T_5581_63; // @[Reg.scala 19:20:@3208.4]
  reg [31:0] _RAND_544;
  wire  _GEN_479; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_480; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_481; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_482; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_483; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_484; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_485; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_486; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_487; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_488; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_489; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_490; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_491; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_492; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_493; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_494; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_495; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_496; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_497; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_498; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_499; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_500; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_501; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_502; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_503; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_504; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_505; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_506; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_507; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_508; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_509; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_510; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_511; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_512; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_513; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_514; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_515; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_516; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_517; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_518; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_519; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_520; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_521; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_522; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_523; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_524; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_525; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_526; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_527; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_528; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_529; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_530; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_531; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_532; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_533; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_534; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_535; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_536; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_537; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_538; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_539; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_540; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_541; // @[Reg.scala 20:19:@3209.4]
  wire  _GEN_542; // @[Reg.scala 20:19:@3209.4]
  reg [7:0] _T_5779; // @[Reg.scala 11:16:@3339.4]
  reg [31:0] _RAND_545;
  reg [7:0] _T_5781; // @[Reg.scala 11:16:@3344.4]
  reg [31:0] _RAND_546;
  reg [7:0] _T_5783; // @[Reg.scala 11:16:@3349.4]
  reg [31:0] _RAND_547;
  reg [7:0] _T_5785; // @[Reg.scala 11:16:@3354.4]
  reg [31:0] _RAND_548;
  reg [7:0] _T_5787; // @[Reg.scala 11:16:@3359.4]
  reg [31:0] _RAND_549;
  reg [7:0] _T_5789; // @[Reg.scala 11:16:@3364.4]
  reg [31:0] _RAND_550;
  reg [7:0] _T_5791; // @[Reg.scala 11:16:@3369.4]
  reg [31:0] _RAND_551;
  reg [7:0] _T_5793; // @[Reg.scala 11:16:@3374.4]
  reg [31:0] _RAND_552;
  reg [7:0] _T_5795; // @[Reg.scala 11:16:@3379.4]
  reg [31:0] _RAND_553;
  reg [7:0] _T_5797; // @[Reg.scala 11:16:@3384.4]
  reg [31:0] _RAND_554;
  reg [7:0] _T_5799; // @[Reg.scala 11:16:@3389.4]
  reg [31:0] _RAND_555;
  reg [7:0] _T_5801; // @[Reg.scala 11:16:@3394.4]
  reg [31:0] _RAND_556;
  reg [7:0] _T_5803; // @[Reg.scala 11:16:@3399.4]
  reg [31:0] _RAND_557;
  reg [7:0] _T_5805; // @[Reg.scala 11:16:@3404.4]
  reg [31:0] _RAND_558;
  reg [7:0] _T_5807; // @[Reg.scala 11:16:@3409.4]
  reg [31:0] _RAND_559;
  reg [7:0] _T_5809; // @[Reg.scala 11:16:@3414.4]
  reg [31:0] _RAND_560;
  reg [7:0] _T_5811; // @[Reg.scala 11:16:@3419.4]
  reg [31:0] _RAND_561;
  reg [7:0] _T_5813; // @[Reg.scala 11:16:@3424.4]
  reg [31:0] _RAND_562;
  reg [7:0] _T_5815; // @[Reg.scala 11:16:@3429.4]
  reg [31:0] _RAND_563;
  reg [7:0] _T_5817; // @[Reg.scala 11:16:@3434.4]
  reg [31:0] _RAND_564;
  reg [7:0] _T_5819; // @[Reg.scala 11:16:@3439.4]
  reg [31:0] _RAND_565;
  reg [7:0] _T_5821; // @[Reg.scala 11:16:@3444.4]
  reg [31:0] _RAND_566;
  reg [7:0] _T_5823; // @[Reg.scala 11:16:@3449.4]
  reg [31:0] _RAND_567;
  reg [7:0] _T_5825; // @[Reg.scala 11:16:@3454.4]
  reg [31:0] _RAND_568;
  reg [7:0] _T_5827; // @[Reg.scala 11:16:@3459.4]
  reg [31:0] _RAND_569;
  reg [7:0] _T_5829; // @[Reg.scala 11:16:@3464.4]
  reg [31:0] _RAND_570;
  reg [7:0] _T_5831; // @[Reg.scala 11:16:@3469.4]
  reg [31:0] _RAND_571;
  reg [7:0] _T_5833; // @[Reg.scala 11:16:@3474.4]
  reg [31:0] _RAND_572;
  reg [7:0] _T_5835; // @[Reg.scala 11:16:@3479.4]
  reg [31:0] _RAND_573;
  reg [7:0] _T_5837; // @[Reg.scala 11:16:@3484.4]
  reg [31:0] _RAND_574;
  reg [7:0] _T_5839; // @[Reg.scala 11:16:@3489.4]
  reg [31:0] _RAND_575;
  reg [7:0] _T_5841; // @[Reg.scala 11:16:@3494.4]
  reg [31:0] _RAND_576;
  reg [7:0] _T_5843; // @[Reg.scala 11:16:@3499.4]
  reg [31:0] _RAND_577;
  reg [7:0] _T_5845; // @[Reg.scala 11:16:@3504.4]
  reg [31:0] _RAND_578;
  reg [7:0] _T_5847; // @[Reg.scala 11:16:@3509.4]
  reg [31:0] _RAND_579;
  reg [7:0] _T_5849; // @[Reg.scala 11:16:@3514.4]
  reg [31:0] _RAND_580;
  reg [7:0] _T_5851; // @[Reg.scala 11:16:@3519.4]
  reg [31:0] _RAND_581;
  reg [7:0] _T_5853; // @[Reg.scala 11:16:@3524.4]
  reg [31:0] _RAND_582;
  reg [7:0] _T_5855; // @[Reg.scala 11:16:@3529.4]
  reg [31:0] _RAND_583;
  reg [7:0] _T_5857; // @[Reg.scala 11:16:@3534.4]
  reg [31:0] _RAND_584;
  reg [7:0] _T_5859; // @[Reg.scala 11:16:@3539.4]
  reg [31:0] _RAND_585;
  reg [7:0] _T_5861; // @[Reg.scala 11:16:@3544.4]
  reg [31:0] _RAND_586;
  reg [7:0] _T_5863; // @[Reg.scala 11:16:@3549.4]
  reg [31:0] _RAND_587;
  reg [7:0] _T_5865; // @[Reg.scala 11:16:@3554.4]
  reg [31:0] _RAND_588;
  reg [7:0] _T_5867; // @[Reg.scala 11:16:@3559.4]
  reg [31:0] _RAND_589;
  reg [7:0] _T_5869; // @[Reg.scala 11:16:@3564.4]
  reg [31:0] _RAND_590;
  reg [7:0] _T_5871; // @[Reg.scala 11:16:@3569.4]
  reg [31:0] _RAND_591;
  reg [7:0] _T_5873; // @[Reg.scala 11:16:@3574.4]
  reg [31:0] _RAND_592;
  reg [7:0] _T_5875; // @[Reg.scala 11:16:@3579.4]
  reg [31:0] _RAND_593;
  reg [7:0] _T_5877; // @[Reg.scala 11:16:@3584.4]
  reg [31:0] _RAND_594;
  reg [7:0] _T_5879; // @[Reg.scala 11:16:@3589.4]
  reg [31:0] _RAND_595;
  reg [7:0] _T_5881; // @[Reg.scala 11:16:@3594.4]
  reg [31:0] _RAND_596;
  reg [7:0] _T_5883; // @[Reg.scala 11:16:@3599.4]
  reg [31:0] _RAND_597;
  reg [7:0] _T_5885; // @[Reg.scala 11:16:@3604.4]
  reg [31:0] _RAND_598;
  reg [7:0] _T_5887; // @[Reg.scala 11:16:@3609.4]
  reg [31:0] _RAND_599;
  reg [7:0] _T_5889; // @[Reg.scala 11:16:@3614.4]
  reg [31:0] _RAND_600;
  reg [7:0] _T_5891; // @[Reg.scala 11:16:@3619.4]
  reg [31:0] _RAND_601;
  reg [7:0] _T_5893; // @[Reg.scala 11:16:@3624.4]
  reg [31:0] _RAND_602;
  reg [7:0] _T_5895; // @[Reg.scala 11:16:@3629.4]
  reg [31:0] _RAND_603;
  reg [7:0] _T_5897; // @[Reg.scala 11:16:@3634.4]
  reg [31:0] _RAND_604;
  reg [7:0] _T_5899; // @[Reg.scala 11:16:@3639.4]
  reg [31:0] _RAND_605;
  reg [7:0] _T_5901; // @[Reg.scala 11:16:@3644.4]
  reg [31:0] _RAND_606;
  reg [7:0] _T_5903; // @[Reg.scala 11:16:@3649.4]
  reg [31:0] _RAND_607;
  reg [7:0] _T_5905; // @[Reg.scala 11:16:@3654.4]
  reg [31:0] _RAND_608;
  reg [7:0] _T_5907; // @[Reg.scala 11:16:@3659.4]
  reg [31:0] _RAND_609;
  reg [7:0] _T_5909; // @[Reg.scala 11:16:@3664.4]
  reg [31:0] _RAND_610;
  reg [7:0] _T_5911; // @[Reg.scala 11:16:@3669.4]
  reg [31:0] _RAND_611;
  reg [7:0] _T_5913; // @[Reg.scala 11:16:@3674.4]
  reg [31:0] _RAND_612;
  reg [7:0] _T_5915; // @[Reg.scala 11:16:@3679.4]
  reg [31:0] _RAND_613;
  reg [7:0] _T_5917; // @[Reg.scala 11:16:@3684.4]
  reg [31:0] _RAND_614;
  reg [7:0] _T_5919; // @[Reg.scala 11:16:@3689.4]
  reg [31:0] _RAND_615;
  reg [7:0] _T_5921; // @[Reg.scala 11:16:@3694.4]
  reg [31:0] _RAND_616;
  reg [7:0] _T_5923; // @[Reg.scala 11:16:@3699.4]
  reg [31:0] _RAND_617;
  reg [7:0] _T_5925; // @[Reg.scala 11:16:@3704.4]
  reg [31:0] _RAND_618;
  reg [7:0] _T_5927; // @[Reg.scala 11:16:@3709.4]
  reg [31:0] _RAND_619;
  reg [7:0] _T_5929; // @[Reg.scala 11:16:@3714.4]
  reg [31:0] _RAND_620;
  reg [7:0] _T_5931; // @[Reg.scala 11:16:@3719.4]
  reg [31:0] _RAND_621;
  reg [7:0] _T_5933; // @[Reg.scala 11:16:@3724.4]
  reg [31:0] _RAND_622;
  reg [7:0] _T_5935; // @[Reg.scala 11:16:@3729.4]
  reg [31:0] _RAND_623;
  reg [7:0] _T_5937; // @[Reg.scala 11:16:@3734.4]
  reg [31:0] _RAND_624;
  reg [7:0] _T_5939; // @[Reg.scala 11:16:@3739.4]
  reg [31:0] _RAND_625;
  reg [7:0] _T_5941; // @[Reg.scala 11:16:@3744.4]
  reg [31:0] _RAND_626;
  reg [7:0] _T_5943; // @[Reg.scala 11:16:@3749.4]
  reg [31:0] _RAND_627;
  reg [7:0] _T_5945; // @[Reg.scala 11:16:@3754.4]
  reg [31:0] _RAND_628;
  reg [7:0] _T_5947; // @[Reg.scala 11:16:@3759.4]
  reg [31:0] _RAND_629;
  reg [7:0] _T_5949; // @[Reg.scala 11:16:@3764.4]
  reg [31:0] _RAND_630;
  reg [7:0] _T_5951; // @[Reg.scala 11:16:@3769.4]
  reg [31:0] _RAND_631;
  reg [7:0] _T_5953; // @[Reg.scala 11:16:@3774.4]
  reg [31:0] _RAND_632;
  reg [7:0] _T_5955; // @[Reg.scala 11:16:@3779.4]
  reg [31:0] _RAND_633;
  reg [7:0] _T_5957; // @[Reg.scala 11:16:@3784.4]
  reg [31:0] _RAND_634;
  reg [7:0] _T_5959; // @[Reg.scala 11:16:@3789.4]
  reg [31:0] _RAND_635;
  reg [7:0] _T_5961; // @[Reg.scala 11:16:@3794.4]
  reg [31:0] _RAND_636;
  reg [7:0] _T_5963; // @[Reg.scala 11:16:@3799.4]
  reg [31:0] _RAND_637;
  reg [7:0] _T_5965; // @[Reg.scala 11:16:@3804.4]
  reg [31:0] _RAND_638;
  reg [7:0] _T_5967; // @[Reg.scala 11:16:@3809.4]
  reg [31:0] _RAND_639;
  reg [7:0] _T_5969; // @[Reg.scala 11:16:@3814.4]
  reg [31:0] _RAND_640;
  reg [7:0] _T_5971; // @[Reg.scala 11:16:@3819.4]
  reg [31:0] _RAND_641;
  reg [7:0] _T_5973; // @[Reg.scala 11:16:@3824.4]
  reg [31:0] _RAND_642;
  reg [7:0] _T_5975; // @[Reg.scala 11:16:@3829.4]
  reg [31:0] _RAND_643;
  reg [7:0] _T_5977; // @[Reg.scala 11:16:@3834.4]
  reg [31:0] _RAND_644;
  reg [7:0] _T_5979; // @[Reg.scala 11:16:@3839.4]
  reg [31:0] _RAND_645;
  reg [7:0] _T_5981; // @[Reg.scala 11:16:@3844.4]
  reg [31:0] _RAND_646;
  reg [7:0] _T_5983; // @[Reg.scala 11:16:@3849.4]
  reg [31:0] _RAND_647;
  reg [7:0] _T_5985; // @[Reg.scala 11:16:@3854.4]
  reg [31:0] _RAND_648;
  reg [7:0] _T_5987; // @[Reg.scala 11:16:@3859.4]
  reg [31:0] _RAND_649;
  reg [7:0] _T_5989; // @[Reg.scala 11:16:@3864.4]
  reg [31:0] _RAND_650;
  reg [7:0] _T_5991; // @[Reg.scala 11:16:@3869.4]
  reg [31:0] _RAND_651;
  reg [7:0] _T_5993; // @[Reg.scala 11:16:@3874.4]
  reg [31:0] _RAND_652;
  reg [7:0] _T_5995; // @[Reg.scala 11:16:@3879.4]
  reg [31:0] _RAND_653;
  reg [7:0] _T_5997; // @[Reg.scala 11:16:@3884.4]
  reg [31:0] _RAND_654;
  reg [7:0] _T_5999; // @[Reg.scala 11:16:@3889.4]
  reg [31:0] _RAND_655;
  reg [7:0] _T_6001; // @[Reg.scala 11:16:@3894.4]
  reg [31:0] _RAND_656;
  reg [7:0] _T_6003; // @[Reg.scala 11:16:@3899.4]
  reg [31:0] _RAND_657;
  reg [7:0] _T_6005; // @[Reg.scala 11:16:@3904.4]
  reg [31:0] _RAND_658;
  reg [7:0] _T_6007; // @[Reg.scala 11:16:@3909.4]
  reg [31:0] _RAND_659;
  reg [7:0] _T_6009; // @[Reg.scala 11:16:@3914.4]
  reg [31:0] _RAND_660;
  reg [7:0] _T_6011; // @[Reg.scala 11:16:@3919.4]
  reg [31:0] _RAND_661;
  reg [7:0] _T_6013; // @[Reg.scala 11:16:@3924.4]
  reg [31:0] _RAND_662;
  reg [7:0] _T_6015; // @[Reg.scala 11:16:@3929.4]
  reg [31:0] _RAND_663;
  reg [7:0] _T_6017; // @[Reg.scala 11:16:@3934.4]
  reg [31:0] _RAND_664;
  reg [7:0] _T_6019; // @[Reg.scala 11:16:@3939.4]
  reg [31:0] _RAND_665;
  reg [7:0] _T_6021; // @[Reg.scala 11:16:@3944.4]
  reg [31:0] _RAND_666;
  reg [7:0] _T_6023; // @[Reg.scala 11:16:@3949.4]
  reg [31:0] _RAND_667;
  reg [7:0] _T_6025; // @[Reg.scala 11:16:@3954.4]
  reg [31:0] _RAND_668;
  reg [7:0] _T_6027; // @[Reg.scala 11:16:@3959.4]
  reg [31:0] _RAND_669;
  reg [7:0] _T_6029; // @[Reg.scala 11:16:@3964.4]
  reg [31:0] _RAND_670;
  reg [7:0] _T_6031; // @[Reg.scala 11:16:@3969.4]
  reg [31:0] _RAND_671;
  reg [7:0] _T_6033; // @[Reg.scala 11:16:@3974.4]
  reg [31:0] _RAND_672;
  assign _T_623 = io_nvdla_core_rstn == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 73:38:@8.4]
  assign _T_625 = io_sc_state == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 77:31:@9.4]
  assign _T_629 = io_sc_state == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 79:31:@11.4]
  assign _T_633 = io_reg2dp_op_en & _T_625; // @[NV_NVDLA_CSC_dl_for_check.scala 86:32:@14.4]
  assign _T_637 = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 88:35:@16.4]
  assign _T_638 = _T_637 & io_reg2dp_datain_format; // @[NV_NVDLA_CSC_dl_for_check.scala 89:22:@17.4]
  assign _T_643 = 7'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_dl_for_check.scala 96:53:@18.4]
  assign _T_645 = _T_638 ? _T_643 : 7'h8; // @[NV_NVDLA_CSC_dl_for_check.scala 96:24:@19.4]
  assign _T_646 = _T_645[5:3]; // @[NV_NVDLA_CSC_dl_for_check.scala 96:100:@20.4]
  assign _T_648 = _T_638 ? _T_646 : 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 97:22:@21.4]
  assign _T_650 = _T_648 - 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 98:34:@22.4]
  assign _T_651 = $unsigned(_T_650); // @[NV_NVDLA_CSC_dl_for_check.scala 98:34:@23.4]
  assign _T_653 = io_reg2dp_conv_x_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 99:51:@24.4]
  assign _T_654 = io_reg2dp_datain_channel_ext[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 100:62:@25.4]
  assign _T_657 = {_T_653,2'h0}; // @[Cat.scala 30:58:@26.4]
  assign _T_660 = {_T_653,1'h0}; // @[Cat.scala 30:58:@27.4]
  assign _GEN_671 = {{1'd0}, _T_653}; // @[NV_NVDLA_CSC_dl_for_check.scala 102:74:@28.4]
  assign _T_661 = _T_660 + _GEN_671; // @[NV_NVDLA_CSC_dl_for_check.scala 102:74:@28.4]
  assign _T_662 = 2'h2 == _T_654; // @[Mux.scala 46:19:@29.4]
  assign _T_663 = _T_662 ? _T_661 : {{2'd0}, _T_653}; // @[Mux.scala 46:16:@30.4]
  assign _T_664 = 2'h3 == _T_654; // @[Mux.scala 46:19:@31.4]
  assign _T_665 = _T_664 ? _T_657 : _T_663; // @[Mux.scala 46:16:@32.4]
  assign _T_667 = io_reg2dp_weight_channel_ext >= 13'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 104:88:@33.4]
  assign _T_673 = io_reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 104:172:@35.4]
  assign _T_674 = _T_667 ? 6'h3f : _T_673; // @[NV_NVDLA_CSC_dl_for_check.scala 104:58:@36.4]
  assign _T_677 = {_T_665,1'h0}; // @[Cat.scala 30:58:@37.4]
  assign _GEN_672 = {{1'd0}, _T_665}; // @[NV_NVDLA_CSC_dl_for_check.scala 105:81:@38.4]
  assign _T_678 = _T_677 + _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 105:81:@38.4]
  assign _T_679 = _T_677 + _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 105:81:@39.4]
  assign _GEN_673 = {{1'd0}, _T_673}; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@41.4]
  assign _T_681 = _T_679 + _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@41.4]
  assign _T_682 = _T_679 + _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@42.4]
  assign _T_685 = _T_665 + _T_673; // @[NV_NVDLA_CSC_dl_for_check.scala 106:58:@44.4]
  assign _T_686 = _T_665 + _T_673; // @[NV_NVDLA_CSC_dl_for_check.scala 106:58:@45.4]
  assign _T_687 = 2'h1 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@46.4]
  assign _T_688 = _T_687 ? _T_686 : _T_674; // @[Mux.scala 46:16:@47.4]
  assign _T_689 = 2'h2 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@48.4]
  assign _T_690 = _T_689 ? _T_682 : {{1'd0}, _T_688}; // @[Mux.scala 46:16:@49.4]
  assign _T_693 = _T_673 + 6'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 107:80:@51.4]
  assign _T_696 = {_T_665,2'h0}; // @[Cat.scala 30:58:@52.4]
  assign _T_701 = _T_687 ? _T_677 : {{1'd0}, _T_665}; // @[Mux.scala 46:16:@55.4]
  assign _T_703 = _T_689 ? _T_696 : {{1'd0}, _T_701}; // @[Mux.scala 46:16:@57.4]
  assign _T_705 = {_T_665,6'h0}; // @[Cat.scala 30:58:@58.4]
  assign _T_707 = io_reg2dp_conv_y_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 117:52:@59.4]
  assign _T_710 = io_reg2dp_x_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 118:60:@60.4]
  assign _T_711 = _T_638 ? 6'h1 : _T_710; // @[NV_NVDLA_CSC_dl_for_check.scala 118:21:@61.4]
  assign _T_714 = io_reg2dp_y_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 119:60:@62.4]
  assign _T_715 = _T_638 ? 6'h1 : _T_714; // @[NV_NVDLA_CSC_dl_for_check.scala 119:21:@63.4]
  assign _T_797 = io_reg2dp_entries + 14'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 135:43:@87.4]
  assign _T_799 = _T_797 * 15'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 136:41:@89.4]
  assign _T_800 = _T_799[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 136:56:@90.4]
  assign _T_801 = 6'h1 * _T_715; // @[NV_NVDLA_CSC_dl_for_check.scala 138:37:@91.4]
  assign _GEN_674 = {{9'd0}, _T_725}; // @[NV_NVDLA_CSC_dl_for_check.scala 139:34:@92.4]
  assign _T_802 = _T_746 * _GEN_674; // @[NV_NVDLA_CSC_dl_for_check.scala 139:34:@92.4]
  assign _T_803 = _T_802[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 139:47:@93.4]
  assign _GEN_675 = {{1'd0}, _T_739}; // @[NV_NVDLA_CSC_dl_for_check.scala 140:34:@94.4]
  assign _T_804 = _T_746 * _GEN_675; // @[NV_NVDLA_CSC_dl_for_check.scala 140:34:@94.4]
  assign _T_805 = _T_804[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 140:51:@95.4]
  assign _T_807 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 141:41:@96.4]
  assign _T_808 = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 141:41:@97.4]
  assign _T_810 = io_reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 142:77:@98.4]
  assign _GEN_676 = {{1'd0}, io_reg2dp_rls_slices}; // @[NV_NVDLA_CSC_dl_for_check.scala 142:113:@99.4]
  assign _T_811 = io_reg2dp_datain_height_ext - _GEN_676; // @[NV_NVDLA_CSC_dl_for_check.scala 142:113:@99.4]
  assign _T_812 = $unsigned(_T_811); // @[NV_NVDLA_CSC_dl_for_check.scala 142:113:@100.4]
  assign _T_813 = io_reg2dp_skip_data_rls ? _T_810 : _T_812; // @[NV_NVDLA_CSC_dl_for_check.scala 142:23:@101.4]
  assign _T_814 = _T_718 ? _T_732 : _T_795; // @[NV_NVDLA_CSC_dl_for_check.scala 143:24:@102.4]
  assign _GEN_677 = {{1'd0}, _T_814}; // @[NV_NVDLA_CSC_dl_for_check.scala 144:38:@103.4]
  assign _T_815 = _T_753 * _GEN_677; // @[NV_NVDLA_CSC_dl_for_check.scala 144:38:@103.4]
  assign _T_816 = _T_815[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 144:54:@104.4]
  assign _T_1041 = _T_638 ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@175.6]
  assign _T_1043 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 193:38:@177.6]
  assign _T_1044 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 193:38:@178.6]
  assign _T_1046 = io_reg2dp_datain_width_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 194:48:@180.6]
  assign _T_1052 = io_reg2dp_weight_channel_ext[12:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 197:93:@185.6]
  assign _T_1053 = {4'h0,_T_1052}; // @[Cat.scala 30:58:@186.6]
  assign _T_1057 = {1'h0,io_reg2dp_entries}; // @[Cat.scala 30:58:@219.6]
  assign _GEN_1 = _T_633 ? _T_1041 : _T_834; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_2 = _T_633 ? _T_1044 : _T_841; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_3 = _T_633 ? _T_1046 : _T_848; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_4 = _T_633 ? io_reg2dp_datain_width_ext : _T_855; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_5 = _T_633 ? io_reg2dp_datain_height_ext : _T_862; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_6 = _T_633 ? _T_1053 : _T_869; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_7 = _T_633 ? _T_646 : _T_872; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_8 = _T_633 ? _T_646 : _T_875; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_10 = _T_633 ? _T_646 : _T_881; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_11 = _T_633 ? _T_646 : _T_884; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_12 = _T_633 ? _T_646 : _T_887; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_13 = _T_633 ? _T_646 : _T_890; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_15 = _T_633 ? _T_646 : _T_896; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_16 = _T_633 ? _T_646 : _T_899; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_18 = _T_633 ? _T_646 : _T_905; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_19 = _T_633 ? _T_648 : _T_908; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_20 = _T_633 ? _T_648 : _T_911; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_21 = _T_633 ? _T_653 : _T_918; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_22 = _T_633 ? _T_707 : _T_925; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_24 = _T_633 ? 6'h1 : _T_725; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_25 = _T_633 ? 5'h0 : _T_935; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_26 = _T_633 ? _T_690 : _T_942; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_27 = _T_633 ? _T_693 : _T_949; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_28 = _T_633 ? _T_703 : _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_29 = _T_633 ? {{1'd0}, _T_665} : _T_963; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_30 = _T_633 ? _T_705 : _T_970; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_31 = _T_633 ? _T_711 : _T_977; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_32 = _T_633 ? _T_715 : _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_33 = _T_633 ? io_reg2dp_pad_value : _T_991; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_34 = _T_633 ? _T_797 : _T_746; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_35 = _T_633 ? _T_800 : _T_753; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_36 = _T_633 ? _T_1057 : _T_998; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_37 = _T_633 ? {{2'd0}, _T_801} : _T_739; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_38 = _T_633 ? {{2'd0}, _T_808} : _T_732; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_39 = _T_633 ? _T_813 : _T_795; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_40 = _T_633 ? io_reg2dp_dataout_width : _T_760; // @[NV_NVDLA_CSC_dl_for_check.scala 190:15:@171.4]
  assign _GEN_43 = _T_718 ? _T_803 : _T_781; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  assign _GEN_44 = _T_718 ? _T_805 : _T_788; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  assign _GEN_45 = _T_718 ? _T_746 : _T_1005; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  assign _GEN_46 = _T_718 ? _T_746 : _T_1012; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  assign _GEN_47 = _T_718 ? _T_816 : _T_774; // @[NV_NVDLA_CSC_dl_for_check.scala 235:18:@232.4]
  assign _GEN_48 = _T_629 ? _T_795 : _T_1019; // @[NV_NVDLA_CSC_dl_for_check.scala 242:17:@239.4]
  assign _GEN_49 = _T_629 ? _T_816 : _T_1026; // @[NV_NVDLA_CSC_dl_for_check.scala 242:17:@239.4]
  assign _T_1159 = _T_1019 != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 306:37:@314.4]
  assign _T_1160 = io_sg2dl_reuse_rls & _T_1159; // @[NV_NVDLA_CSC_dl_for_check.scala 306:23:@315.4]
  assign _T_2244 = _T_881[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 896:32:@1229.4]
  assign _T_2245 = _T_2244 & _T_2220; // @[NV_NVDLA_CSC_dl_for_check.scala 896:36:@1230.4]
  assign _T_2246 = _T_881[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 897:35:@1231.4]
  assign _T_2247 = _T_2246 & _T_2214; // @[NV_NVDLA_CSC_dl_for_check.scala 897:39:@1232.4]
  assign _T_2248 = _T_2245 | _T_2247; // @[NV_NVDLA_CSC_dl_for_check.scala 896:57:@1233.4]
  assign _T_2249 = _T_881[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 898:35:@1234.4]
  assign _T_2250 = _T_2249 & _T_2211; // @[NV_NVDLA_CSC_dl_for_check.scala 898:39:@1235.4]
  assign _T_2251 = _T_2248 | _T_2250; // @[NV_NVDLA_CSC_dl_for_check.scala 897:60:@1236.4]
  assign _T_2252 = _T_884[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 905:42:@1238.4]
  assign _T_2256 = _T_2252 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1240.4]
  assign _T_2257 = _T_2256 & _T_2234; // @[NV_NVDLA_CSC_dl_for_check.scala 905:47:@1241.4]
  assign _T_2258 = _T_884[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 906:42:@1242.4]
  assign _T_2262 = _T_2258 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1244.4]
  assign _T_2263 = _T_2262 & _T_2228; // @[NV_NVDLA_CSC_dl_for_check.scala 906:47:@1245.4]
  assign _T_2264 = _T_2257 | _T_2263; // @[NV_NVDLA_CSC_dl_for_check.scala 905:66:@1246.4]
  assign _T_2265 = _T_884[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 907:42:@1247.4]
  assign _T_2269 = _T_2265 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1249.4]
  assign _T_2270 = _T_2269 & _T_2225; // @[NV_NVDLA_CSC_dl_for_check.scala 907:47:@1250.4]
  assign _T_2271 = _T_2264 | _T_2270; // @[NV_NVDLA_CSC_dl_for_check.scala 906:66:@1251.4]
  assign _T_2290 = _T_2271[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 931:26:@1270.4]
  assign _T_1157 = _T_2251 & _T_2290; // @[NV_NVDLA_CSC_dl_for_check.scala 303:29:@313.4]
  assign _T_1162 = _T_732 != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 306:66:@316.4]
  assign _T_1163 = _T_1157 & _T_1162; // @[NV_NVDLA_CSC_dl_for_check.scala 306:53:@317.4]
  assign _T_1164 = _T_1160 | _T_1163; // @[NV_NVDLA_CSC_dl_for_check.scala 306:42:@318.4]
  assign _T_1165 = _T_1157 ? _T_732 : _T_1019; // @[NV_NVDLA_CSC_dl_for_check.scala 307:28:@320.4]
  assign _T_1166 = _T_1157 ? _T_774 : _T_1026; // @[NV_NVDLA_CSC_dl_for_check.scala 308:29:@322.4]
  assign _T_1097 = _T_1164 ? _T_1166 : 15'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 275:28:@262.4]
  assign _T_1105 = _T_1079 + _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 280:37:@269.4]
  assign _T_1106 = _T_1079 + _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 280:37:@270.4]
  assign _T_1112 = {_T_841,9'h0}; // @[Cat.scala 30:58:@272.4]
  assign _GEN_678 = {{1'd0}, _T_1112}; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@273.4]
  assign _T_1113 = _T_1106 - _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@273.4]
  assign _T_1114 = $unsigned(_T_1113); // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@274.4]
  assign _T_1115 = _T_1114[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 281:46:@275.4]
  assign _T_1122 = _T_1106 >= _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 282:45:@278.4]
  assign _T_1124 = _T_1122 ? _T_1115 : _T_1106; // @[NV_NVDLA_CSC_dl_for_check.scala 283:83:@279.4]
  assign _T_1125 = io_sc2cdma_dat_pending_req ? 15'h0 : _T_1124; // @[NV_NVDLA_CSC_dl_for_check.scala 283:25:@280.4]
  assign _T_1151 = _T_1164 | io_sc2cdma_dat_pending_req; // @[NV_NVDLA_CSC_dl_for_check.scala 294:13:@303.4]
  assign _GEN_52 = _T_1151 ? _T_1125 : _T_1079; // @[NV_NVDLA_CSC_dl_for_check.scala 294:25:@304.4]
  assign _GEN_54 = _T_1164 ? _T_1165 : _T_1172; // @[Reg.scala 20:19:@328.4]
  assign _GEN_55 = _T_1164 ? _T_1166 : _T_1175; // @[Reg.scala 20:19:@333.4]
  assign _T_1225 = {{30'd0}, _T_1192}; // @[NV_NVDLA_CSC_dl_for_check.scala 343:19:@376.4 NV_NVDLA_CSC_dl_for_check.scala 347:12:@382.4]
  assign _GEN_61 = _T_1192 ? _T_1225 : _T_1228; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@384.4]
  assign _GEN_62 = _T_1214 ? _T_1228 : _T_1231; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@388.4]
  assign _GEN_63 = _T_1217 ? _T_1231 : _T_1234; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@392.4]
  assign _GEN_64 = _T_1220 ? _T_1234 : _T_1237; // @[NV_NVDLA_CSC_dl_for_check.scala 351:23:@396.4]
  assign _T_1238 = _T_872[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 356:30:@399.4]
  assign _T_1239 = _T_1238 & _T_1214; // @[NV_NVDLA_CSC_dl_for_check.scala 356:34:@400.4]
  assign _T_1240 = _T_872[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 357:30:@401.4]
  assign _T_1241 = _T_1240 & _T_1220; // @[NV_NVDLA_CSC_dl_for_check.scala 357:34:@402.4]
  assign _T_1242 = _T_1239 | _T_1241; // @[NV_NVDLA_CSC_dl_for_check.scala 356:50:@403.4]
  assign _T_1243 = _T_872[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 358:30:@404.4]
  assign _T_1244 = _T_1243 & _T_1223; // @[NV_NVDLA_CSC_dl_for_check.scala 358:34:@405.4]
  assign _T_1245 = _T_1242 | _T_1244; // @[NV_NVDLA_CSC_dl_for_check.scala 357:50:@406.4]
  assign _T_1246 = _T_875[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 360:37:@407.4]
  assign _T_1250 = _T_1246 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@409.4]
  assign _T_1251 = _T_1250 & _T_1228; // @[NV_NVDLA_CSC_dl_for_check.scala 360:42:@410.4]
  assign _T_1252 = _T_875[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 361:37:@411.4]
  assign _T_1256 = _T_1252 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@413.4]
  assign _T_1257 = _T_1256 & _T_1234; // @[NV_NVDLA_CSC_dl_for_check.scala 361:42:@414.4]
  assign _T_1258 = _T_1251 | _T_1257; // @[NV_NVDLA_CSC_dl_for_check.scala 360:56:@415.4]
  assign _T_1259 = _T_875[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 362:37:@416.4]
  assign _T_1263 = _T_1259 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@418.4]
  assign _T_1264 = _T_1263 & _T_1237; // @[NV_NVDLA_CSC_dl_for_check.scala 362:42:@419.4]
  assign _T_1265 = _T_1258 | _T_1264; // @[NV_NVDLA_CSC_dl_for_check.scala 361:56:@420.4]
  assign _T_1266 = _T_1265[4:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 365:24:@421.4]
  assign _T_1267 = _T_1265[9:5]; // @[NV_NVDLA_CSC_dl_for_check.scala 366:24:@422.4]
  assign _T_1268 = _T_1265[16:10]; // @[NV_NVDLA_CSC_dl_for_check.scala 367:28:@423.4]
  assign _T_1269 = _T_1265[23:17]; // @[NV_NVDLA_CSC_dl_for_check.scala 368:29:@424.4]
  assign _T_1270 = _T_1265[25:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 369:25:@425.4]
  assign _T_1271 = _T_1265[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 370:25:@426.4]
  assign _T_1272 = _T_1265[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 371:27:@427.4]
  assign _T_1273 = _T_1265[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 372:25:@428.4]
  assign _T_1274 = _T_1265[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 373:25:@429.4]
  assign _T_1275 = _T_1265[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 374:27:@430.4]
  assign _T_1286 = _T_1282 + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 383:24:@434.4]
  assign _T_1287 = _T_1282 + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 383:24:@435.4]
  assign _T_1290 = _T_1282 == _T_935; // @[NV_NVDLA_CSC_dl_for_check.scala 385:27:@439.4]
  assign _T_1288 = _T_1290 ? 5'h0 : _T_1287; // @[NV_NVDLA_CSC_dl_for_check.scala 382:17:@436.4]
  assign _T_1289 = _T_633 ? 5'h0 : _T_1288; // @[NV_NVDLA_CSC_dl_for_check.scala 381:17:@437.4]
  assign _T_1297 = _T_1293 + 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 391:31:@443.4]
  assign _T_1298 = _T_1293 + 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 391:31:@444.4]
  assign _GEN_682 = {{1'd0}, _T_1298}; // @[NV_NVDLA_CSC_dl_for_check.scala 392:32:@445.4]
  assign _T_1299 = _GEN_682 == _T_908; // @[NV_NVDLA_CSC_dl_for_check.scala 392:32:@445.4]
  assign _T_1301 = io_reg2dp_y_extension != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 393:61:@447.4]
  assign _T_1349 = _T_1309 != 7'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 426:37:@484.4]
  assign _T_1350 = ~ _T_1349; // @[NV_NVDLA_CSC_dl_for_check.scala 426:24:@485.4]
  assign _T_1352 = _T_1293 != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 426:56:@486.4]
  assign _T_1353 = ~ _T_1352; // @[NV_NVDLA_CSC_dl_for_check.scala 426:44:@487.4]
  assign _T_1354 = _T_1350 & _T_1353; // @[NV_NVDLA_CSC_dl_for_check.scala 426:42:@488.4]
  assign _T_1356 = _T_1282 != 5'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 426:75:@489.4]
  assign _T_1357 = ~ _T_1356; // @[NV_NVDLA_CSC_dl_for_check.scala 426:63:@490.4]
  assign _T_1358 = _T_1354 & _T_1357; // @[NV_NVDLA_CSC_dl_for_check.scala 426:61:@491.4]
  assign _T_1360 = _T_1358 ? 1'h0 : _T_1338; // @[NV_NVDLA_CSC_dl_for_check.scala 426:22:@492.4]
  assign _T_1361 = _T_1245 ? 1'h1 : _T_1360; // @[NV_NVDLA_CSC_dl_for_check.scala 425:22:@493.4]
  assign _T_1302 = _T_1301 & _T_1361; // @[NV_NVDLA_CSC_dl_for_check.scala 393:66:@448.4]
  assign _T_1303 = _T_633 | _T_1302; // @[NV_NVDLA_CSC_dl_for_check.scala 393:33:@449.4]
  assign _T_1304 = _T_633 | _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 395:31:@451.6]
  assign _T_1306 = _T_1304 ? 2'h0 : _T_1298; // @[NV_NVDLA_CSC_dl_for_check.scala 395:21:@452.6]
  assign _GEN_65 = _T_1303 ? _T_1306 : _T_1293; // @[NV_NVDLA_CSC_dl_for_check.scala 394:23:@450.4]
  assign _T_1315 = _T_1309 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 403:33:@458.4]
  assign _T_1316 = _T_1309 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 403:33:@459.4]
  assign _T_1317 = _T_1316 == _T_1269; // @[NV_NVDLA_CSC_dl_for_check.scala 404:51:@460.4]
  assign _T_1318 = _T_1290 & _T_1317; // @[NV_NVDLA_CSC_dl_for_check.scala 404:33:@461.4]
  assign _T_1319 = _T_1318 & _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 405:34:@463.4]
  assign _T_1320 = _T_1361 & _T_1290; // @[NV_NVDLA_CSC_dl_for_check.scala 406:52:@465.4]
  assign _T_1321 = _T_633 | _T_1320; // @[NV_NVDLA_CSC_dl_for_check.scala 406:34:@466.4]
  assign _T_1323 = ~ _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 410:41:@468.6]
  assign _T_1324 = _T_1318 & _T_1323; // @[NV_NVDLA_CSC_dl_for_check.scala 410:39:@469.6]
  assign _T_1327 = _T_1319 ? 7'h0 : _T_1316; // @[NV_NVDLA_CSC_dl_for_check.scala 411:22:@470.6]
  assign _T_1328 = _T_1324 ? 7'h0 : _T_1327; // @[NV_NVDLA_CSC_dl_for_check.scala 410:22:@471.6]
  assign _T_1329 = _T_633 ? 7'h0 : _T_1328; // @[NV_NVDLA_CSC_dl_for_check.scala 409:22:@472.6]
  assign _GEN_66 = _T_1321 ? _T_1329 : _T_1309; // @[NV_NVDLA_CSC_dl_for_check.scala 408:24:@467.4]
  assign _T_1346 = _T_1245 | _T_1332; // @[NV_NVDLA_CSC_dl_for_check.scala 424:27:@482.4]
  assign _T_1341 = _T_1346 & _T_1318; // @[NV_NVDLA_CSC_dl_for_check.scala 421:49:@479.4]
  assign _T_1344 = _T_1245 ? 1'h1 : _T_1332; // @[NV_NVDLA_CSC_dl_for_check.scala 422:32:@480.4]
  assign _T_1345 = _T_1341 ? 1'h0 : _T_1344; // @[NV_NVDLA_CSC_dl_for_check.scala 421:33:@481.4]
  assign _T_1366 = {1'h0,_T_1268}; // @[Cat.scala 30:58:@499.4]
  assign _GEN_67 = _T_1361 ? _T_1366 : _T_1364; // @[NV_NVDLA_CSC_dl_for_check.scala 436:21:@500.4]
  assign _GEN_683 = {{10'd0}, _T_911}; // @[NV_NVDLA_CSC_dl_for_check.scala 446:39:@505.4]
  assign _T_1373 = _T_1369 + _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 446:39:@505.4]
  assign _T_1374 = _T_1369 + _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 446:39:@506.4]
  assign _T_1375 = _T_1290 & _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 447:29:@507.4]
  assign _T_1376 = _T_1369 >= _T_760; // @[NV_NVDLA_CSC_dl_for_check.scala 447:61:@508.4]
  assign _T_1377 = _T_1375 & _T_1376; // @[NV_NVDLA_CSC_dl_for_check.scala 447:44:@509.4]
  assign _T_1380 = ~ _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 450:43:@512.4]
  assign _T_1381 = _T_1319 & _T_1380; // @[NV_NVDLA_CSC_dl_for_check.scala 450:41:@513.4]
  assign _T_1382 = _T_1377 ? {{9'd0}, _T_651} : _T_1374; // @[NV_NVDLA_CSC_dl_for_check.scala 451:26:@514.4]
  assign _T_1383 = _T_1381 ? _T_1372 : _T_1382; // @[NV_NVDLA_CSC_dl_for_check.scala 450:26:@515.4]
  assign _T_1384 = _T_633 ? {{9'd0}, _T_651} : _T_1383; // @[NV_NVDLA_CSC_dl_for_check.scala 449:26:@516.4]
  assign _T_1386 = _T_1320 & _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 452:70:@518.4]
  assign _T_1387 = _T_633 | _T_1386; // @[NV_NVDLA_CSC_dl_for_check.scala 452:37:@519.4]
  assign _T_1388 = _T_1361 & _T_1319; // @[NV_NVDLA_CSC_dl_for_check.scala 453:55:@520.4]
  assign _T_1389 = _T_1388 & _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 453:71:@521.4]
  assign _T_1390 = _T_633 | _T_1389; // @[NV_NVDLA_CSC_dl_for_check.scala 453:37:@522.4]
  assign _GEN_68 = _T_1387 ? _T_1384 : _T_1369; // @[NV_NVDLA_CSC_dl_for_check.scala 455:27:@523.4]
  assign _GEN_69 = _T_1390 ? _T_1384 : _T_1372; // @[NV_NVDLA_CSC_dl_for_check.scala 458:27:@526.4]
  assign _T_1394 = _T_1393 == _T_869; // @[NV_NVDLA_CSC_dl_for_check.scala 465:37:@530.4]
  assign _T_1396 = _T_1388 & _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 466:70:@532.4]
  assign _T_1397 = _T_633 | _T_1396; // @[NV_NVDLA_CSC_dl_for_check.scala 466:36:@533.4]
  assign _T_1401 = _T_1393 + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 471:34:@535.6]
  assign _T_1402 = _T_1393 + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 471:34:@536.6]
  assign _T_1403 = _T_1272 ? 11'h0 : _T_1402; // @[NV_NVDLA_CSC_dl_for_check.scala 470:24:@537.6]
  assign _T_1404 = _T_633 ? 11'h0 : _T_1403; // @[NV_NVDLA_CSC_dl_for_check.scala 469:24:@538.6]
  assign _GEN_70 = _T_1397 ? _T_1404 : _T_1393; // @[NV_NVDLA_CSC_dl_for_check.scala 468:26:@534.4]
  assign _GEN_684 = {{8'd0}, io_reg2dp_pad_left}; // @[NV_NVDLA_CSC_dl_for_check.scala 486:41:@550.4]
  assign _T_1433 = 13'h0 - _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 486:41:@550.4]
  assign _T_1434 = $unsigned(_T_1433); // @[NV_NVDLA_CSC_dl_for_check.scala 486:41:@551.4]
  assign _T_1435 = _T_638 ? 14'h0 : _T_1434; // @[NV_NVDLA_CSC_dl_for_check.scala 485:26:@552.4]
  assign _GEN_685 = {{10'd0}, _T_918}; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@553.4]
  assign _T_1436 = _T_1407 + _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@553.4]
  assign _T_1437 = _T_1407 + _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@554.4]
  assign _T_1440 = _T_1377 ? _T_1435 : _T_1437; // @[NV_NVDLA_CSC_dl_for_check.scala 492:25:@557.4]
  assign _T_1441 = _T_1381 ? _T_1410 : _T_1440; // @[NV_NVDLA_CSC_dl_for_check.scala 491:25:@558.4]
  assign _T_1442 = _T_633 ? _T_1435 : _T_1441; // @[NV_NVDLA_CSC_dl_for_check.scala 490:25:@559.4]
  assign _GEN_686 = {{1'd0}, _T_1266}; // @[NV_NVDLA_CSC_dl_for_check.scala 494:35:@560.4]
  assign _T_1443 = _GEN_686 * _T_977; // @[NV_NVDLA_CSC_dl_for_check.scala 494:35:@560.4]
  assign _GEN_687 = {{3'd0}, _T_1443}; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@561.4]
  assign _T_1444 = _T_1407 + _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@561.4]
  assign _T_1445 = _T_1407 + _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@562.4]
  assign _T_1448 = _T_834[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 496:96:@565.4]
  assign _T_1449 = ~ _T_1448; // @[NV_NVDLA_CSC_dl_for_check.scala 496:86:@566.4]
  assign _T_1450 = _T_1386 & _T_1449; // @[NV_NVDLA_CSC_dl_for_check.scala 496:84:@567.4]
  assign _T_1451 = _T_633 | _T_1450; // @[NV_NVDLA_CSC_dl_for_check.scala 496:36:@568.4]
  assign _T_1454 = _T_834[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 497:99:@571.4]
  assign _T_1455 = ~ _T_1454; // @[NV_NVDLA_CSC_dl_for_check.scala 497:89:@572.4]
  assign _T_1456 = _T_1389 & _T_1455; // @[NV_NVDLA_CSC_dl_for_check.scala 497:87:@573.4]
  assign _T_1457 = _T_633 | _T_1456; // @[NV_NVDLA_CSC_dl_for_check.scala 497:36:@574.4]
  assign _T_1459 = _T_1299 ? _T_956 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 500:26:@575.4]
  assign _T_1462 = _T_673 == 6'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 502:79:@577.4]
  assign _T_1466 = _T_1052 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 503:74:@580.4]
  assign _T_1467 = _T_1052 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 503:74:@581.4]
  assign _T_1468 = _T_1462 ? _T_1052 : _T_1467; // @[NV_NVDLA_CSC_dl_for_check.scala 502:27:@582.4]
  assign _T_1469 = _T_1272 & _T_1319; // @[NV_NVDLA_CSC_dl_for_check.scala 504:37:@583.4]
  assign _T_1471 = _T_1271 & _T_1319; // @[NV_NVDLA_CSC_dl_for_check.scala 505:35:@584.4]
  assign _T_1473 = _T_1422 + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 505:66:@585.4]
  assign _T_1474 = _T_1422 + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 505:66:@586.4]
  assign _T_1475 = _T_1471 ? _T_1474 : _T_1422; // @[NV_NVDLA_CSC_dl_for_check.scala 505:22:@587.4]
  assign _T_1476 = _T_1469 ? 13'h2 : _T_1475; // @[NV_NVDLA_CSC_dl_for_check.scala 504:22:@588.4]
  assign _GEN_688 = {{6'd0}, _T_1468}; // @[NV_NVDLA_CSC_dl_for_check.scala 507:44:@590.4]
  assign _T_1477 = _T_1422 >= _GEN_688; // @[NV_NVDLA_CSC_dl_for_check.scala 507:44:@590.4]
  assign _T_1478 = _T_1319 & _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 511:39:@591.4]
  assign _T_1479 = _T_1478 & _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 511:54:@592.4]
  assign _T_1480 = _T_1479 & _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 511:71:@593.4]
  assign _T_1483 = ~ _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 512:73:@596.4]
  assign _T_1484 = _T_1479 & _T_1483; // @[NV_NVDLA_CSC_dl_for_check.scala 512:71:@597.4]
  assign _GEN_689 = {{4'd0}, _T_970}; // @[NV_NVDLA_CSC_dl_for_check.scala 512:99:@598.4]
  assign _T_1485 = _T_1419 + _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 512:99:@598.4]
  assign _T_1486 = _T_1419 + _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 512:99:@599.4]
  assign _T_1488 = _T_1478 & _T_1477; // @[NV_NVDLA_CSC_dl_for_check.scala 513:54:@601.4]
  assign _GEN_690 = {{9'd0}, _T_949}; // @[NV_NVDLA_CSC_dl_for_check.scala 513:90:@602.4]
  assign _T_1489 = _T_1416 + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 513:90:@602.4]
  assign _T_1490 = _T_1416 + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 513:90:@603.4]
  assign _T_1492 = ~ _T_1477; // @[NV_NVDLA_CSC_dl_for_check.scala 514:56:@605.4]
  assign _T_1493 = _T_1478 & _T_1492; // @[NV_NVDLA_CSC_dl_for_check.scala 514:54:@606.4]
  assign _T_1495 = _T_1416 + 16'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 514:91:@607.4]
  assign _T_1496 = _T_1416 + 16'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 514:91:@608.4]
  assign _T_1497 = ~ _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 515:41:@609.4]
  assign _T_1498 = _T_1319 & _T_1497; // @[NV_NVDLA_CSC_dl_for_check.scala 515:39:@610.4]
  assign _GEN_691 = {{8'd0}, _T_1459}; // @[NV_NVDLA_CSC_dl_for_check.scala 515:81:@611.4]
  assign _T_1499 = _T_1413 + _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 515:81:@611.4]
  assign _T_1500 = _T_1413 + _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 515:81:@612.4]
  assign _T_1501 = _T_1498 ? _T_1416 : _T_1500; // @[NV_NVDLA_CSC_dl_for_check.scala 515:24:@613.4]
  assign _T_1502 = _T_1493 ? _T_1496 : _T_1501; // @[NV_NVDLA_CSC_dl_for_check.scala 514:24:@614.4]
  assign _T_1503 = _T_1488 ? _T_1490 : _T_1502; // @[NV_NVDLA_CSC_dl_for_check.scala 513:24:@615.4]
  assign _T_1504 = _T_1484 ? _T_1486 : _T_1503; // @[NV_NVDLA_CSC_dl_for_check.scala 512:24:@616.4]
  assign _T_1505 = _T_1480 ? {{9'd0}, _T_942} : _T_1504; // @[NV_NVDLA_CSC_dl_for_check.scala 511:24:@617.4]
  assign _T_1506 = _T_718 ? {{9'd0}, _T_942} : _T_1505; // @[NV_NVDLA_CSC_dl_for_check.scala 510:24:@618.4]
  assign _T_1512 = _T_1413[15:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 517:68:@620.4]
  assign _T_1513 = {5'h0,_T_1512}; // @[Cat.scala 30:58:@621.4]
  assign _T_1524 = _T_834[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 520:68:@632.4]
  assign _T_1525 = _T_1361 & _T_1524; // @[NV_NVDLA_CSC_dl_for_check.scala 520:57:@633.4]
  assign _T_1526 = _T_1525 & _T_1319; // @[NV_NVDLA_CSC_dl_for_check.scala 520:72:@634.4]
  assign _T_1527 = _T_1526 & _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 520:88:@635.4]
  assign _T_1528 = _T_1527 & _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 520:103:@636.4]
  assign _T_1529 = _T_718 | _T_1528; // @[NV_NVDLA_CSC_dl_for_check.scala 520:39:@637.4]
  assign _T_1531 = _T_1448 & _T_1245; // @[NV_NVDLA_CSC_dl_for_check.scala 522:42:@639.4]
  assign _T_1534 = _T_1427 ? 1'h0 : _T_1430; // @[NV_NVDLA_CSC_dl_for_check.scala 522:74:@640.4]
  assign _T_1535 = _T_1531 ? 1'h1 : _T_1534; // @[NV_NVDLA_CSC_dl_for_check.scala 522:28:@641.4]
  assign _T_1537 = _T_1448 & _T_1299; // @[NV_NVDLA_CSC_dl_for_check.scala 523:36:@643.4]
  assign _T_1538 = _T_1535 | _T_1430; // @[NV_NVDLA_CSC_dl_for_check.scala 523:72:@644.4]
  assign _T_1539 = _T_1537 & _T_1538; // @[NV_NVDLA_CSC_dl_for_check.scala 523:51:@645.4]
  assign _GEN_71 = _T_1451 ? _T_1442 : _T_1407; // @[NV_NVDLA_CSC_dl_for_check.scala 525:26:@646.4]
  assign _GEN_72 = _T_1451 ? _T_1506 : _T_1413; // @[NV_NVDLA_CSC_dl_for_check.scala 525:26:@646.4]
  assign _GEN_73 = _T_1457 ? _T_1442 : _T_1410; // @[NV_NVDLA_CSC_dl_for_check.scala 529:26:@650.4]
  assign _GEN_74 = _T_1457 ? _T_1506 : _T_1416; // @[NV_NVDLA_CSC_dl_for_check.scala 529:26:@650.4]
  assign _GEN_75 = _T_1529 ? _T_1506 : _T_1419; // @[NV_NVDLA_CSC_dl_for_check.scala 533:26:@654.4]
  assign _GEN_692 = {{9'd0}, io_reg2dp_pad_top}; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@659.4]
  assign _T_1547 = 14'h0 - _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@659.4]
  assign _T_1548 = $unsigned(_T_1547); // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@660.4]
  assign _T_1549 = _T_1548[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 542:41:@661.4]
  assign _GEN_693 = {{10'd0}, _T_925}; // @[NV_NVDLA_CSC_dl_for_check.scala 543:37:@662.4]
  assign _T_1550 = _T_1542 + _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 543:37:@662.4]
  assign _T_1551 = _T_1542 + _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 543:37:@663.4]
  assign _T_1552 = _T_1319 & _T_1273; // @[NV_NVDLA_CSC_dl_for_check.scala 544:52:@664.4]
  assign _T_1553 = _T_633 | _T_1552; // @[NV_NVDLA_CSC_dl_for_check.scala 544:35:@665.4]
  assign _T_1556 = _T_1377 ? _T_1551 : _T_1542; // @[NV_NVDLA_CSC_dl_for_check.scala 546:25:@668.4]
  assign _T_1557 = _T_1381 ? _T_1545 : _T_1556; // @[NV_NVDLA_CSC_dl_for_check.scala 545:25:@669.4]
  assign _T_1558 = _T_1553 ? _T_1549 : _T_1557; // @[NV_NVDLA_CSC_dl_for_check.scala 544:25:@670.4]
  assign _T_1561 = _T_1381 | _T_1377; // @[NV_NVDLA_CSC_dl_for_check.scala 547:91:@673.4]
  assign _T_1562 = _T_1361 & _T_1561; // @[NV_NVDLA_CSC_dl_for_check.scala 547:54:@674.4]
  assign _T_1563 = _T_633 | _T_1562; // @[NV_NVDLA_CSC_dl_for_check.scala 547:36:@675.4]
  assign _GEN_694 = {{1'd0}, _T_1267}; // @[NV_NVDLA_CSC_dl_for_check.scala 549:35:@679.4]
  assign _T_1567 = _GEN_694 * _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 549:35:@679.4]
  assign _GEN_695 = {{3'd0}, _T_1567}; // @[NV_NVDLA_CSC_dl_for_check.scala 550:33:@680.4]
  assign _T_1568 = _T_1542 + _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 550:33:@680.4]
  assign _T_1569 = _T_1542 + _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 550:33:@681.4]
  assign _GEN_696 = {{12'd0}, _T_1293}; // @[NV_NVDLA_CSC_dl_for_check.scala 550:51:@682.4]
  assign _T_1570 = _T_1569 + _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 550:51:@682.4]
  assign _T_1571 = _T_1569 + _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 550:51:@683.4]
  assign _GEN_76 = _T_1563 ? _T_1558 : _T_1542; // @[NV_NVDLA_CSC_dl_for_check.scala 552:26:@684.4]
  assign _GEN_77 = _T_1390 ? _T_1558 : _T_1545; // @[NV_NVDLA_CSC_dl_for_check.scala 553:26:@687.4]
  assign _T_1572 = _T_1445[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 556:39:@690.4]
  assign _GEN_697 = {{1'd0}, _T_855}; // @[NV_NVDLA_CSC_dl_for_check.scala 556:59:@691.4]
  assign _T_1573 = _T_1445 > _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 556:59:@691.4]
  assign _T_1574 = _T_1572 | _T_1573; // @[NV_NVDLA_CSC_dl_for_check.scala 556:44:@692.4]
  assign _T_1575 = _T_1571[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 556:92:@693.4]
  assign _T_1576 = _T_1574 | _T_1575; // @[NV_NVDLA_CSC_dl_for_check.scala 556:78:@694.4]
  assign _GEN_698 = {{1'd0}, _T_862}; // @[NV_NVDLA_CSC_dl_for_check.scala 556:112:@695.4]
  assign _T_1577 = _T_1571 > _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 556:112:@695.4]
  assign _T_1578 = _T_1576 | _T_1577; // @[NV_NVDLA_CSC_dl_for_check.scala 556:97:@696.4]
  assign _T_1591 = _T_1575 | _T_1577; // @[NV_NVDLA_CSC_dl_for_check.scala 559:42:@706.4]
  assign _T_1701 = _T_834[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 644:33:@792.4]
  assign _T_1702 = ~ _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 645:24:@793.4]
  assign _T_1704 = _T_1445[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 645:77:@794.4]
  assign _T_1705 = {2'h0,_T_1704}; // @[Cat.scala 30:58:@795.4]
  assign _T_1707 = _T_1366 > 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 646:38:@796.4]
  assign _T_1712 = _T_1445[12:1]; // @[NV_NVDLA_CSC_dl_for_check.scala 647:54:@799.4]
  assign _T_1713 = {3'h0,_T_1712}; // @[Cat.scala 30:58:@800.4]
  assign _T_1714 = _T_1707 ? _T_1705 : _T_1713; // @[NV_NVDLA_CSC_dl_for_check.scala 646:23:@801.4]
  assign _T_1715 = _T_1702 ? _T_1705 : _T_1714; // @[NV_NVDLA_CSC_dl_for_check.scala 645:23:@802.4]
  assign _T_1716 = _T_1701 ? _T_1513 : _T_1715; // @[NV_NVDLA_CSC_dl_for_check.scala 644:23:@803.4]
  assign _T_1717 = _T_1716[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 656:24:@805.4]
  assign _T_1594 = _T_1717[13:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 563:32:@708.4]
  assign _GEN_700 = {{3'd0}, _T_1594}; // @[NV_NVDLA_CSC_dl_for_check.scala 563:40:@709.4]
  assign _T_1595 = _GEN_700 > _T_998; // @[NV_NVDLA_CSC_dl_for_check.scala 563:40:@709.4]
  assign _T_1596 = _T_834[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 564:34:@710.4]
  assign _T_1597 = _T_1596 ? _T_1591 : _T_1578; // @[NV_NVDLA_CSC_dl_for_check.scala 564:24:@711.4]
  assign _T_1598 = _T_834[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 565:29:@712.4]
  assign _T_1599 = _T_1598 & _T_1595; // @[NV_NVDLA_CSC_dl_for_check.scala 565:33:@713.4]
  assign _T_1600 = ~ _T_1597; // @[NV_NVDLA_CSC_dl_for_check.scala 566:39:@714.4]
  assign _T_1601 = _T_1361 & _T_1600; // @[NV_NVDLA_CSC_dl_for_check.scala 566:37:@715.4]
  assign _T_1602 = ~ _T_1599; // @[NV_NVDLA_CSC_dl_for_check.scala 566:56:@716.4]
  assign _T_1603 = _T_1601 & _T_1602; // @[NV_NVDLA_CSC_dl_for_check.scala 566:54:@717.4]
  assign _T_1604 = _T_834[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 569:37:@718.4]
  assign _T_1605 = ~ _T_1604; // @[NV_NVDLA_CSC_dl_for_check.scala 569:27:@719.4]
  assign _T_1606 = _T_1393[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 569:54:@720.4]
  assign _T_1607 = _T_1605 ? _T_1606 : _T_1271; // @[NV_NVDLA_CSC_dl_for_check.scala 569:26:@721.4]
  assign _T_1608 = _T_1445[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 570:35:@722.4]
  assign _T_1610 = _T_1293 == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 571:55:@723.4]
  assign _T_1611 = _T_1361 & _T_1610; // @[NV_NVDLA_CSC_dl_for_check.scala 571:42:@724.4]
  assign _T_1612 = _T_1318 & _T_1346; // @[NV_NVDLA_CSC_dl_for_check.scala 574:42:@726.4]
  assign _T_1616 = {_T_1274,_T_1272,_T_1612,_T_1245,_T_1282}; // @[Cat.scala 30:58:@730.4]
  assign _T_1647 = _T_1275 & _T_1318; // @[NV_NVDLA_CSC_dl_for_check.scala 601:38:@750.6]
  assign _T_1648 = _T_1647 & _T_1346; // @[NV_NVDLA_CSC_dl_for_check.scala 601:56:@751.6]
  assign _GEN_78 = _T_1361 ? _T_1608 : _T_1622; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_79 = _T_1361 ? _T_1293 : _T_1625; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_80 = _T_1361 ? _T_1607 : _T_1628; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_81 = _T_1361 ? _T_1394 : _T_1631; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_82 = _T_1361 ? _T_1361 : _T_1634; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_83 = _T_1361 ? _T_1270 : _T_1637; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_84 = _T_1361 ? _T_1616 : _T_1643; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_85 = _T_1361 ? _T_1648 : _T_1646; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_86 = _T_1361 ? _T_1535 : _T_1430; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_87 = _T_1361 ? _T_1539 : _T_1427; // @[NV_NVDLA_CSC_dl_for_check.scala 593:21:@742.4]
  assign _GEN_88 = _T_1611 ? _T_1245 : _T_1640; // @[NV_NVDLA_CSC_dl_for_check.scala 605:26:@756.4]
  assign _T_1670 = _T_834[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 622:32:@766.4]
  assign _T_1671 = ~ _T_1670; // @[NV_NVDLA_CSC_dl_for_check.scala 622:22:@767.4]
  assign _T_1672 = _T_848[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 622:49:@768.4]
  assign _T_1674 = _T_1671 ? _T_1672 : 12'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 622:21:@769.4]
  assign _T_1676 = _T_1319 & _T_1272; // @[NV_NVDLA_CSC_dl_for_check.scala 624:34:@770.4]
  assign _GEN_701 = {{1'd0}, _T_1674}; // @[NV_NVDLA_CSC_dl_for_check.scala 624:64:@771.4]
  assign _T_1678 = _T_1651 + _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 624:64:@771.4]
  assign _T_1679 = _T_1651 + _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 624:64:@772.4]
  assign _T_1680 = _T_1676 ? 13'h0 : _T_1679; // @[NV_NVDLA_CSC_dl_for_check.scala 624:19:@773.4]
  assign _T_1681 = _T_633 ? 13'h0 : _T_1680; // @[NV_NVDLA_CSC_dl_for_check.scala 623:19:@774.4]
  assign _T_1685 = _T_1651 != _T_1654; // @[NV_NVDLA_CSC_dl_for_check.scala 626:31:@778.4]
  assign _GEN_702 = {{2'd0}, _T_781}; // @[NV_NVDLA_CSC_dl_for_check.scala 629:32:@779.4]
  assign _T_1686 = _T_1542 * _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 629:32:@779.4]
  assign _T_1687 = _T_1686[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 629:50:@780.4]
  assign _GEN_703 = {{7'd0}, _T_1267}; // @[NV_NVDLA_CSC_dl_for_check.scala 630:31:@781.4]
  assign _T_1688 = _GEN_703 * _T_788; // @[NV_NVDLA_CSC_dl_for_check.scala 630:31:@781.4]
  assign _T_1689 = _T_1688[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 630:49:@782.4]
  assign _GEN_704 = {{10'd0}, _T_1282}; // @[NV_NVDLA_CSC_dl_for_check.scala 631:29:@783.4]
  assign _T_1690 = _GEN_704 * _T_1005; // @[NV_NVDLA_CSC_dl_for_check.scala 631:29:@783.4]
  assign _T_1691 = _T_1690[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 631:47:@784.4]
  assign _GEN_705 = {{13'd0}, _T_1293}; // @[NV_NVDLA_CSC_dl_for_check.scala 632:47:@785.4]
  assign _T_1693 = _GEN_705 * _T_1012; // @[NV_NVDLA_CSC_dl_for_check.scala 632:47:@785.4]
  assign _T_1694 = _T_633 ? 17'h0 : _T_1693; // @[NV_NVDLA_CSC_dl_for_check.scala 632:21:@786.4]
  assign _T_1695 = _T_1694[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 632:65:@787.4]
  assign _T_1696 = _T_834[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 633:45:@788.4]
  assign _T_1697 = _T_633 | _T_1696; // @[NV_NVDLA_CSC_dl_for_check.scala 633:34:@789.4]
  assign _T_1698 = {_T_1697,_T_1361}; // @[Cat.scala 30:58:@790.4]
  assign _GEN_89 = _T_1397 ? _T_1681 : _T_1651; // @[NV_NVDLA_CSC_dl_for_check.scala 660:20:@807.4]
  assign _GEN_90 = _T_1685 ? _T_1651 : _T_1654; // @[NV_NVDLA_CSC_dl_for_check.scala 663:23:@810.4]
  assign _T_1718 = _T_1698[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 666:19:@813.4]
  assign _GEN_91 = _T_1718 ? _T_1687 : _T_1657; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@814.4]
  assign _GEN_92 = _T_1718 ? _T_1689 : _T_1660; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@814.4]
  assign _GEN_93 = _T_1718 ? _T_1691 : _T_1663; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@814.4]
  assign _T_1719 = _T_1698[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 671:19:@819.4]
  assign _GEN_94 = _T_1719 ? _T_1695 : _T_1666; // @[NV_NVDLA_CSC_dl_for_check.scala 671:23:@820.4]
  assign _GEN_95 = _T_1361 ? _T_1717 : {{1'd0}, _T_1669}; // @[NV_NVDLA_CSC_dl_for_check.scala 674:20:@823.4]
  assign _T_1825 = _T_1657 + _T_1660; // @[NV_NVDLA_CSC_dl_for_check.scala 698:29:@851.4]
  assign _T_1826 = _T_1657 + _T_1660; // @[NV_NVDLA_CSC_dl_for_check.scala 698:29:@852.4]
  assign _T_1827 = _T_1826 + _T_1663; // @[NV_NVDLA_CSC_dl_for_check.scala 698:43:@853.4]
  assign _T_1828 = _T_1826 + _T_1663; // @[NV_NVDLA_CSC_dl_for_check.scala 698:43:@854.4]
  assign _T_1829 = _T_1828 + _T_1666; // @[NV_NVDLA_CSC_dl_for_check.scala 698:57:@855.4]
  assign _T_1830 = _T_1828 + _T_1666; // @[NV_NVDLA_CSC_dl_for_check.scala 698:57:@856.4]
  assign _GEN_706 = {{2'd0}, _T_1654}; // @[NV_NVDLA_CSC_dl_for_check.scala 699:40:@857.4]
  assign _T_1831 = _T_1079 + _GEN_706; // @[NV_NVDLA_CSC_dl_for_check.scala 699:40:@857.4]
  assign _T_1832 = _T_1079 + _GEN_706; // @[NV_NVDLA_CSC_dl_for_check.scala 699:40:@858.4]
  assign _GEN_707 = {{2'd0}, _T_1830}; // @[NV_NVDLA_CSC_dl_for_check.scala 699:52:@859.4]
  assign _T_1833 = _T_1832 + _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 699:52:@859.4]
  assign _T_1834 = _T_1832 + _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 699:52:@860.4]
  assign _GEN_708 = {{2'd0}, _T_1669}; // @[NV_NVDLA_CSC_dl_for_check.scala 699:64:@861.4]
  assign _T_1835 = _T_1834 + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 699:64:@861.4]
  assign _T_1836 = _T_1834 + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 699:64:@862.4]
  assign _T_1843 = _T_1836 >= _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 700:45:@865.4]
  assign _T_1850 = _T_1836 - _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 701:42:@868.4]
  assign _T_1851 = $unsigned(_T_1850); // @[NV_NVDLA_CSC_dl_for_check.scala 701:42:@869.4]
  assign _T_1852 = _T_1851[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 701:42:@870.4]
  assign _T_1853 = _T_633 | _T_1634; // @[NV_NVDLA_CSC_dl_for_check.scala 702:35:@871.4]
  assign _T_1859 = _T_1843 ? _T_1852 : _T_1836; // @[NV_NVDLA_CSC_dl_for_check.scala 703:25:@873.4]
  assign _T_1860 = _T_1853 ? 15'h1fff : _T_1859; // @[NV_NVDLA_CSC_dl_for_check.scala 702:25:@874.4]
  assign _T_1884 = 2'h3 == _T_1625; // @[Mux.scala 46:19:@884.4]
  assign _T_1885 = _T_1884 ? _T_1762_3 : 13'h0; // @[Mux.scala 46:16:@885.4]
  assign _T_1886 = 2'h2 == _T_1625; // @[Mux.scala 46:19:@886.4]
  assign _T_1887 = _T_1886 ? _T_1762_2 : _T_1885; // @[Mux.scala 46:16:@887.4]
  assign _T_1888 = 2'h1 == _T_1625; // @[Mux.scala 46:19:@888.4]
  assign _T_1889 = _T_1888 ? _T_1762_1 : _T_1887; // @[Mux.scala 46:16:@889.4]
  assign _T_1890 = 2'h0 == _T_1625; // @[Mux.scala 46:19:@890.4]
  assign _T_1891 = _T_1890 ? _T_1762_0 : _T_1889; // @[Mux.scala 46:16:@891.4]
  assign _GEN_712 = {{2'd0}, _T_1891}; // @[NV_NVDLA_CSC_dl_for_check.scala 710:65:@892.4]
  assign _T_1892 = _GEN_712 != _T_1860; // @[NV_NVDLA_CSC_dl_for_check.scala 710:65:@892.4]
  assign _T_1893 = _T_1892 | _T_1430; // @[NV_NVDLA_CSC_dl_for_check.scala 710:85:@893.4]
  assign _T_1894 = _T_1619 & _T_1893; // @[NV_NVDLA_CSC_dl_for_check.scala 710:43:@894.4]
  assign _T_1895 = _T_1619 | _T_1634; // @[NV_NVDLA_CSC_dl_for_check.scala 712:38:@895.4]
  assign _T_1897 = _T_1625 == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@896.4]
  assign _T_1898 = _T_1895 & _T_1897; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@897.4]
  assign _T_1899 = _T_633 | _T_1898; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@898.4]
  assign _T_1902 = _T_1625 == 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@900.4]
  assign _T_1903 = _T_1895 & _T_1902; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@901.4]
  assign _T_1904 = _T_633 | _T_1903; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@902.4]
  assign _T_1907 = _T_1625 == 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@904.4]
  assign _T_1908 = _T_1895 & _T_1907; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@905.4]
  assign _T_1909 = _T_633 | _T_1908; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@906.4]
  assign _T_1912 = _T_1625 == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 712:78:@908.4]
  assign _T_1913 = _T_1895 & _T_1912; // @[NV_NVDLA_CSC_dl_for_check.scala 712:58:@909.4]
  assign _T_1914 = _T_633 | _T_1913; // @[NV_NVDLA_CSC_dl_for_check.scala 712:17:@910.4]
  assign _GEN_96 = _T_1899 ? _T_1860 : {{2'd0}, _T_1762_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@916.4]
  assign _GEN_97 = _T_1904 ? _T_1860 : {{2'd0}, _T_1762_1}; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@919.4]
  assign _GEN_98 = _T_1909 ? _T_1860 : {{2'd0}, _T_1762_2}; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@922.4]
  assign _GEN_99 = _T_1914 ? _T_1860 : {{2'd0}, _T_1762_3}; // @[NV_NVDLA_CSC_dl_for_check.scala 719:35:@925.4]
  assign _T_1925 = _T_633 | _T_1894; // @[NV_NVDLA_CSC_dl_for_check.scala 725:14:@929.4]
  assign _GEN_100 = _T_1925 ? _T_1860 : _T_1788; // @[NV_NVDLA_CSC_dl_for_check.scala 725:34:@930.4]
  assign _GEN_101 = _T_1338 ? _T_1622 : _T_1797; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_102 = _T_1338 ? _T_1625 : _T_1800; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_103 = _T_1338 ? _T_1628 : _T_1803; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_104 = _T_1338 ? _T_1631 : _T_1806; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_105 = _T_1338 ? _T_1364 : _T_1809; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_106 = _T_1338 ? _T_1634 : _T_1812; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_107 = _T_1338 ? _T_1637 : _T_1815; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_108 = _T_1338 ? _T_1640 : _T_1818; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_109 = _T_1338 ? _T_1646 : _T_1821; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _GEN_110 = _T_1338 ? _T_1643 : {{8'd0}, _T_1338}; // @[NV_NVDLA_CSC_dl_for_check.scala 732:24:@937.4]
  assign _T_1935 = {1'h0,_T_1806,_T_1803,_T_1800,_T_1797}; // @[Cat.scala 30:58:@957.4]
  assign _T_1941 = {_T_1824,_T_1821,_T_1818,_T_1812,_T_1815,_T_1809,_T_1935}; // @[Cat.scala 30:58:@963.4]
  assign _GEN_111 = _T_1791 ? _T_1941 : _T_1966; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1005.4]
  assign _GEN_114 = _T_1946 ? _T_1966 : _T_1969; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1014.4]
  assign _GEN_117 = _T_1949 ? _T_1969 : _T_1972; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1023.4]
  assign _GEN_120 = _T_1952 ? _T_1972 : _T_1975; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1032.4]
  assign _GEN_123 = _T_1955 ? _T_1975 : _T_1978; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1041.4]
  assign _GEN_126 = _T_1958 ? _T_1978 : _T_1981; // @[NV_NVDLA_CSC_dl_for_check.scala 777:33:@1050.4]
  assign _T_2042 = _T_1981[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 794:41:@1058.4]
  assign _T_2043 = _T_1981[3:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 795:41:@1059.4]
  assign _T_2044 = _T_1981[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 796:41:@1060.4]
  assign _T_2045 = _T_1981[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 797:42:@1061.4]
  assign _T_2046 = _T_1981[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 798:41:@1062.4]
  assign _T_2047 = _T_1981[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 799:45:@1063.4]
  assign _T_2050 = _T_1981[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 802:39:@1066.4]
  assign _T_2051 = _T_1981[28:20]; // @[NV_NVDLA_CSC_dl_for_check.scala 803:40:@1067.4]
  assign _T_2108 = _T_834[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 833:69:@1095.4]
  assign _T_2109 = _T_2108 & io_sc2buf_dat_rd_data_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 833:74:@1096.4]
  assign _T_2110 = ~ _T_2054; // @[NV_NVDLA_CSC_dl_for_check.scala 833:90:@1097.4]
  assign _T_2111 = _T_2109 & _T_2110; // @[NV_NVDLA_CSC_dl_for_check.scala 833:88:@1098.4]
  assign _T_2151 = io_sc2buf_dat_rd_data_valid ? 1'h0 : _T_2054; // @[NV_NVDLA_CSC_dl_for_check.scala 848:22:@1132.4]
  assign _T_2165 = io_sc2buf_dat_rd_data_valid ? _T_2054 : _T_2066; // @[NV_NVDLA_CSC_dl_for_check.scala 852:48:@1143.4]
  assign _T_2166 = _T_2111 ? 1'h0 : _T_2165; // @[NV_NVDLA_CSC_dl_for_check.scala 852:22:@1144.4]
  assign _T_2243 = {_T_2051,_T_2050,_T_2047,_T_2046,1'h0,_T_2045,_T_2044,_T_2043,_T_2042}; // @[Cat.scala 30:58:@1211.4]
  assign _GEN_137 = _T_1961 ? _T_2243 : _T_2225; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1214.4]
  assign _GEN_138 = _T_2211 ? _T_2225 : _T_2228; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1218.4]
  assign _GEN_139 = _T_2214 ? _T_2228 : _T_2231; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1222.4]
  assign _GEN_140 = _T_2217 ? _T_2231 : _T_2234; // @[NV_NVDLA_CSC_dl_for_check.scala 891:28:@1226.4]
  assign _T_2272 = _T_2225[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 909:39:@1252.4]
  assign _T_2273 = _T_2228[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 910:39:@1253.4]
  assign _T_2274 = _T_2231[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 911:39:@1254.4]
  assign _T_2275 = _T_2234[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 912:39:@1255.4]
  assign _T_2276 = _T_2225[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 914:38:@1256.4]
  assign _T_2277 = _T_2228[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 915:38:@1257.4]
  assign _T_2278 = _T_2231[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 916:38:@1258.4]
  assign _T_2279 = _T_2234[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 917:38:@1259.4]
  assign _T_2280 = _T_2276[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 919:44:@1260.4]
  assign _T_2281 = _T_2277[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 920:44:@1261.4]
  assign _T_2282 = _T_2278[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 921:44:@1262.4]
  assign _T_2283 = _T_2279[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 922:44:@1263.4]
  assign _T_2284 = _T_2271[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 925:31:@1264.4]
  assign _T_2288 = _T_2271[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 929:31:@1268.4]
  assign _T_2289 = _T_2271[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 930:35:@1269.4]
  assign _T_2299 = io_sc2buf_dat_rd_data_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 941:29:@1278.4]
  assign _T_2310 = _T_963 > 7'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 946:50:@1282.4]
  assign _GEN_713 = {{1'd0}, _T_963}; // @[NV_NVDLA_CSC_dl_for_check.scala 946:111:@1283.4]
  assign _T_2312 = _T_2185 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 946:111:@1283.4]
  assign _T_2313 = _T_2185 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 946:111:@1284.4]
  assign _T_2314 = _T_2313 - _T_2299; // @[NV_NVDLA_CSC_dl_for_check.scala 946:133:@1285.4]
  assign _T_2315 = $unsigned(_T_2314); // @[NV_NVDLA_CSC_dl_for_check.scala 946:133:@1286.4]
  assign _T_2316 = _T_2315[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 946:133:@1287.4]
  assign _T_2317 = _T_2310 ? 8'h40 : _T_2316; // @[NV_NVDLA_CSC_dl_for_check.scala 946:29:@1288.4]
  assign _T_2321 = _T_2188 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 947:111:@1290.4]
  assign _T_2322 = _T_2188 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 947:111:@1291.4]
  assign _T_2323 = _T_2322 - 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 947:133:@1292.4]
  assign _T_2324 = $unsigned(_T_2323); // @[NV_NVDLA_CSC_dl_for_check.scala 947:133:@1293.4]
  assign _T_2325 = _T_2324[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 947:133:@1294.4]
  assign _T_2326 = _T_2310 ? 8'h40 : _T_2325; // @[NV_NVDLA_CSC_dl_for_check.scala 947:29:@1295.4]
  assign _T_2330 = _T_2191 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 948:111:@1297.4]
  assign _T_2331 = _T_2191 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 948:111:@1298.4]
  assign _T_2332 = _T_2331 - 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 948:133:@1299.4]
  assign _T_2333 = $unsigned(_T_2332); // @[NV_NVDLA_CSC_dl_for_check.scala 948:133:@1300.4]
  assign _T_2334 = _T_2333[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 948:133:@1301.4]
  assign _T_2335 = _T_2310 ? 8'h40 : _T_2334; // @[NV_NVDLA_CSC_dl_for_check.scala 948:29:@1302.4]
  assign _T_2339 = _T_2194 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 949:111:@1304.4]
  assign _T_2340 = _T_2194 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 949:111:@1305.4]
  assign _T_2341 = _T_2340 - 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 949:133:@1306.4]
  assign _T_2342 = $unsigned(_T_2341); // @[NV_NVDLA_CSC_dl_for_check.scala 949:133:@1307.4]
  assign _T_2343 = _T_2342[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 949:133:@1308.4]
  assign _T_2344 = _T_2310 ? 8'h40 : _T_2343; // @[NV_NVDLA_CSC_dl_for_check.scala 949:29:@1309.4]
  assign _T_2346 = ~ _T_2272; // @[NV_NVDLA_CSC_dl_for_check.scala 958:52:@1310.4]
  assign _T_2347 = _T_2280 & _T_2346; // @[NV_NVDLA_CSC_dl_for_check.scala 958:50:@1311.4]
  assign _T_2348 = _T_2280 & _T_2272; // @[NV_NVDLA_CSC_dl_for_check.scala 959:50:@1312.4]
  assign _T_2353 = _T_2348 ? 8'h40 : _T_2317; // @[NV_NVDLA_CSC_dl_for_check.scala 959:27:@1315.4]
  assign _T_2354 = _T_2347 ? _T_2197 : _T_2353; // @[NV_NVDLA_CSC_dl_for_check.scala 958:27:@1316.4]
  assign _T_2355 = _T_633 ? 8'h40 : _T_2354; // @[NV_NVDLA_CSC_dl_for_check.scala 957:27:@1317.4]
  assign _T_2357 = ~ _T_2273; // @[NV_NVDLA_CSC_dl_for_check.scala 963:52:@1318.4]
  assign _T_2358 = _T_2281 & _T_2357; // @[NV_NVDLA_CSC_dl_for_check.scala 963:50:@1319.4]
  assign _T_2359 = _T_2281 & _T_2273; // @[NV_NVDLA_CSC_dl_for_check.scala 964:50:@1320.4]
  assign _T_2364 = _T_2359 ? 8'h40 : _T_2326; // @[NV_NVDLA_CSC_dl_for_check.scala 964:27:@1323.4]
  assign _T_2365 = _T_2358 ? _T_2200 : _T_2364; // @[NV_NVDLA_CSC_dl_for_check.scala 963:27:@1324.4]
  assign _T_2366 = _T_633 ? 8'h40 : _T_2365; // @[NV_NVDLA_CSC_dl_for_check.scala 962:27:@1325.4]
  assign _T_2368 = ~ _T_2274; // @[NV_NVDLA_CSC_dl_for_check.scala 968:52:@1326.4]
  assign _T_2369 = _T_2282 & _T_2368; // @[NV_NVDLA_CSC_dl_for_check.scala 968:50:@1327.4]
  assign _T_2370 = _T_2282 & _T_2274; // @[NV_NVDLA_CSC_dl_for_check.scala 969:50:@1328.4]
  assign _T_2375 = _T_2370 ? 8'h40 : _T_2335; // @[NV_NVDLA_CSC_dl_for_check.scala 969:27:@1331.4]
  assign _T_2376 = _T_2369 ? _T_2203 : _T_2375; // @[NV_NVDLA_CSC_dl_for_check.scala 968:27:@1332.4]
  assign _T_2377 = _T_633 ? 8'h40 : _T_2376; // @[NV_NVDLA_CSC_dl_for_check.scala 967:27:@1333.4]
  assign _T_2379 = ~ _T_2275; // @[NV_NVDLA_CSC_dl_for_check.scala 973:52:@1334.4]
  assign _T_2380 = _T_2283 & _T_2379; // @[NV_NVDLA_CSC_dl_for_check.scala 973:50:@1335.4]
  assign _T_2381 = _T_2283 & _T_2275; // @[NV_NVDLA_CSC_dl_for_check.scala 974:50:@1336.4]
  assign _T_2386 = _T_2381 ? 8'h40 : _T_2344; // @[NV_NVDLA_CSC_dl_for_check.scala 974:27:@1339.4]
  assign _T_2387 = _T_2380 ? _T_2206 : _T_2386; // @[NV_NVDLA_CSC_dl_for_check.scala 973:27:@1340.4]
  assign _T_2388 = _T_633 ? 8'h40 : _T_2387; // @[NV_NVDLA_CSC_dl_for_check.scala 972:27:@1341.4]
  assign _T_2389 = _T_834[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 978:46:@1342.4]
  assign _T_2390 = _T_2389 & _T_2211; // @[NV_NVDLA_CSC_dl_for_check.scala 978:51:@1343.4]
  assign _T_2391 = _T_633 | _T_2390; // @[NV_NVDLA_CSC_dl_for_check.scala 978:34:@1344.4]
  assign _T_2392 = _T_834[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 979:46:@1345.4]
  assign _T_2393 = _T_2392 & _T_2214; // @[NV_NVDLA_CSC_dl_for_check.scala 979:51:@1346.4]
  assign _T_2395 = _T_887 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 979:87:@1347.4]
  assign _T_2396 = _T_2393 & _T_2395; // @[NV_NVDLA_CSC_dl_for_check.scala 979:69:@1348.4]
  assign _T_2397 = _T_633 | _T_2396; // @[NV_NVDLA_CSC_dl_for_check.scala 979:34:@1349.4]
  assign _T_2398 = _T_834[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 980:46:@1350.4]
  assign _T_2399 = _T_2398 & _T_2217; // @[NV_NVDLA_CSC_dl_for_check.scala 980:51:@1351.4]
  assign _T_2401 = _T_887 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 980:87:@1352.4]
  assign _T_2402 = _T_2399 & _T_2401; // @[NV_NVDLA_CSC_dl_for_check.scala 980:69:@1353.4]
  assign _T_2403 = _T_633 | _T_2402; // @[NV_NVDLA_CSC_dl_for_check.scala 980:34:@1354.4]
  assign _T_2404 = _T_834[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 981:46:@1355.4]
  assign _T_2405 = _T_2404 & _T_2220; // @[NV_NVDLA_CSC_dl_for_check.scala 981:51:@1356.4]
  assign _T_2408 = _T_2405 & _T_2401; // @[NV_NVDLA_CSC_dl_for_check.scala 981:69:@1358.4]
  assign _T_2409 = _T_633 | _T_2408; // @[NV_NVDLA_CSC_dl_for_check.scala 981:34:@1359.4]
  assign _T_2410 = _T_834[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 983:50:@1360.4]
  assign _T_2411 = _T_2410 & _T_2211; // @[NV_NVDLA_CSC_dl_for_check.scala 983:55:@1361.4]
  assign _T_2412 = _T_2411 & _T_2280; // @[NV_NVDLA_CSC_dl_for_check.scala 983:73:@1362.4]
  assign _T_2413 = _T_2412 & _T_2272; // @[NV_NVDLA_CSC_dl_for_check.scala 983:97:@1363.4]
  assign _T_2414 = _T_633 | _T_2413; // @[NV_NVDLA_CSC_dl_for_check.scala 983:38:@1364.4]
  assign _T_2415 = _T_834[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 984:50:@1365.4]
  assign _T_2416 = _T_2415 & _T_2214; // @[NV_NVDLA_CSC_dl_for_check.scala 984:55:@1366.4]
  assign _T_2417 = _T_2416 & _T_2281; // @[NV_NVDLA_CSC_dl_for_check.scala 984:73:@1367.4]
  assign _T_2418 = _T_2417 & _T_2273; // @[NV_NVDLA_CSC_dl_for_check.scala 984:97:@1368.4]
  assign _T_2420 = _T_890 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 984:138:@1369.4]
  assign _T_2421 = _T_2418 & _T_2420; // @[NV_NVDLA_CSC_dl_for_check.scala 984:120:@1370.4]
  assign _T_2422 = _T_633 | _T_2421; // @[NV_NVDLA_CSC_dl_for_check.scala 984:38:@1371.4]
  assign _T_2423 = _T_834[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 985:50:@1372.4]
  assign _T_2424 = _T_2423 & _T_2217; // @[NV_NVDLA_CSC_dl_for_check.scala 985:55:@1373.4]
  assign _T_2425 = _T_2424 & _T_2282; // @[NV_NVDLA_CSC_dl_for_check.scala 985:73:@1374.4]
  assign _T_2426 = _T_2425 & _T_2274; // @[NV_NVDLA_CSC_dl_for_check.scala 985:97:@1375.4]
  assign _T_2428 = _T_890 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 985:138:@1376.4]
  assign _T_2429 = _T_2426 & _T_2428; // @[NV_NVDLA_CSC_dl_for_check.scala 985:120:@1377.4]
  assign _T_2430 = _T_633 | _T_2429; // @[NV_NVDLA_CSC_dl_for_check.scala 985:38:@1378.4]
  assign _T_2431 = _T_834[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 986:50:@1379.4]
  assign _T_2432 = _T_2431 & _T_2220; // @[NV_NVDLA_CSC_dl_for_check.scala 986:55:@1380.4]
  assign _T_2433 = _T_2432 & _T_2283; // @[NV_NVDLA_CSC_dl_for_check.scala 986:73:@1381.4]
  assign _T_2434 = _T_2433 & _T_2275; // @[NV_NVDLA_CSC_dl_for_check.scala 986:97:@1382.4]
  assign _T_2437 = _T_2434 & _T_2428; // @[NV_NVDLA_CSC_dl_for_check.scala 986:120:@1384.4]
  assign _T_2438 = _T_633 | _T_2437; // @[NV_NVDLA_CSC_dl_for_check.scala 986:38:@1385.4]
  assign _GEN_141 = _T_2391 ? _T_2355 : _T_2185; // @[NV_NVDLA_CSC_dl_for_check.scala 988:24:@1386.4]
  assign _GEN_142 = _T_2397 ? _T_2366 : _T_2188; // @[NV_NVDLA_CSC_dl_for_check.scala 989:24:@1389.4]
  assign _GEN_143 = _T_2403 ? _T_2377 : _T_2191; // @[NV_NVDLA_CSC_dl_for_check.scala 990:24:@1392.4]
  assign _GEN_144 = _T_2409 ? _T_2388 : _T_2194; // @[NV_NVDLA_CSC_dl_for_check.scala 991:24:@1395.4]
  assign _GEN_145 = _T_2414 ? _T_2355 : _T_2197; // @[NV_NVDLA_CSC_dl_for_check.scala 992:28:@1398.4]
  assign _GEN_146 = _T_2422 ? _T_2366 : _T_2200; // @[NV_NVDLA_CSC_dl_for_check.scala 993:28:@1401.4]
  assign _GEN_147 = _T_2430 ? _T_2377 : _T_2203; // @[NV_NVDLA_CSC_dl_for_check.scala 994:28:@1404.4]
  assign _GEN_148 = _T_2438 ? _T_2388 : _T_2206; // @[NV_NVDLA_CSC_dl_for_check.scala 995:28:@1407.4]
  assign _T_2439 = _T_991[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1004:55:@1410.4]
  assign _T_2442 = {_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439}; // @[Cat.scala 30:58:@1413.4]
  assign _T_2443 = {_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2442}; // @[Cat.scala 30:58:@1414.4]
  assign _T_2444 = {_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2439,_T_2442,_T_2443}; // @[Cat.scala 30:58:@1415.4]
  assign _T_2445 = {_T_2444,_T_2444}; // @[Cat.scala 30:58:@1416.4]
  assign _T_2446 = _T_2054 ? _T_2445 : _T_2077; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:23:@1417.4]
  assign _T_2450 = _T_2066 ? _T_2445 : _T_2085; // @[NV_NVDLA_CSC_dl_for_check.scala 1011:23:@1421.4]
  assign _T_2456 = _T_834[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1024:37:@1426.4]
  assign _T_2459 = _T_2288 <= 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:43:@1427.4]
  assign _T_2460 = _T_2284[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:87:@1428.4]
  assign _T_2462 = _T_2460 == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:91:@1429.4]
  assign _T_2463 = _T_2459 & _T_2462; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:72:@1430.4]
  assign _T_2465 = _T_2446[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:171:@1431.4]
  assign _T_2466 = {256'h0,_T_2465}; // @[Cat.scala 30:58:@1432.4]
  assign _T_2472 = _T_2459 & _T_2460; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:72:@1436.4]
  assign _T_2474 = _T_2446[511:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:171:@1437.4]
  assign _T_2475 = {256'h0,_T_2474}; // @[Cat.scala 30:58:@1438.4]
  assign _T_2476 = _T_2472 ? _T_2475 : _T_2446; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:27:@1439.4]
  assign _T_2477 = _T_2463 ? _T_2466 : _T_2476; // @[NV_NVDLA_CSC_dl_for_check.scala 1025:27:@1440.4]
  assign _T_2478 = _T_2456 ? 512'h0 : _T_2477; // @[NV_NVDLA_CSC_dl_for_check.scala 1024:27:@1441.4]
  assign _T_2549 = _T_2478[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1444.4]
  assign _T_2550 = _T_2478[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1446.4]
  assign _T_2551 = _T_2478[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1448.4]
  assign _T_2552 = _T_2478[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1450.4]
  assign _T_2553 = _T_2478[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1452.4]
  assign _T_2554 = _T_2478[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1454.4]
  assign _T_2555 = _T_2478[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1456.4]
  assign _T_2556 = _T_2478[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1458.4]
  assign _T_2557 = _T_2478[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1460.4]
  assign _T_2558 = _T_2478[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1462.4]
  assign _T_2559 = _T_2478[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1464.4]
  assign _T_2560 = _T_2478[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1466.4]
  assign _T_2561 = _T_2478[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1468.4]
  assign _T_2562 = _T_2478[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1470.4]
  assign _T_2563 = _T_2478[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1472.4]
  assign _T_2564 = _T_2478[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1474.4]
  assign _T_2565 = _T_2478[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1476.4]
  assign _T_2566 = _T_2478[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1478.4]
  assign _T_2567 = _T_2478[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1480.4]
  assign _T_2568 = _T_2478[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1482.4]
  assign _T_2569 = _T_2478[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1484.4]
  assign _T_2570 = _T_2478[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1486.4]
  assign _T_2571 = _T_2478[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1488.4]
  assign _T_2572 = _T_2478[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1490.4]
  assign _T_2573 = _T_2478[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1492.4]
  assign _T_2574 = _T_2478[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1494.4]
  assign _T_2575 = _T_2478[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1496.4]
  assign _T_2576 = _T_2478[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1498.4]
  assign _T_2577 = _T_2478[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1500.4]
  assign _T_2578 = _T_2478[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1502.4]
  assign _T_2579 = _T_2478[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1504.4]
  assign _T_2580 = _T_2478[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1506.4]
  assign _T_2581 = _T_2478[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1508.4]
  assign _T_2582 = _T_2478[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1510.4]
  assign _T_2583 = _T_2478[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1512.4]
  assign _T_2584 = _T_2478[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1514.4]
  assign _T_2585 = _T_2478[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1516.4]
  assign _T_2586 = _T_2478[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1518.4]
  assign _T_2587 = _T_2478[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1520.4]
  assign _T_2588 = _T_2478[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1522.4]
  assign _T_2589 = _T_2478[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1524.4]
  assign _T_2590 = _T_2478[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1526.4]
  assign _T_2591 = _T_2478[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1528.4]
  assign _T_2592 = _T_2478[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1530.4]
  assign _T_2593 = _T_2478[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1532.4]
  assign _T_2594 = _T_2478[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1534.4]
  assign _T_2595 = _T_2478[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1536.4]
  assign _T_2596 = _T_2478[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1538.4]
  assign _T_2597 = _T_2478[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1540.4]
  assign _T_2598 = _T_2478[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1542.4]
  assign _T_2599 = _T_2478[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1544.4]
  assign _T_2600 = _T_2478[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1546.4]
  assign _T_2601 = _T_2478[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1548.4]
  assign _T_2602 = _T_2478[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1550.4]
  assign _T_2603 = _T_2478[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1552.4]
  assign _T_2604 = _T_2478[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1554.4]
  assign _T_2605 = _T_2478[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1556.4]
  assign _T_2606 = _T_2478[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1558.4]
  assign _T_2607 = _T_2478[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1560.4]
  assign _T_2608 = _T_2478[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1562.4]
  assign _T_2609 = _T_2478[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1564.4]
  assign _T_2610 = _T_2478[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1566.4]
  assign _T_2611 = _T_2478[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1568.4]
  assign _T_2612 = _T_2478[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1042:39:@1570.4]
  assign _T_2625 = _T_834[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1055:39:@1578.4]
  assign _T_2626 = ~ _T_2625; // @[NV_NVDLA_CSC_dl_for_check.scala 1055:29:@1579.4]
  assign _T_2628 = {_T_2446,_T_2450}; // @[Cat.scala 30:58:@1580.4]
  assign _T_2629 = _T_2626 ? 1024'h0 : _T_2628; // @[NV_NVDLA_CSC_dl_for_check.scala 1055:28:@1581.4]
  assign _T_2630 = _T_834[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1056:39:@1582.4]
  assign _T_2631 = ~ _T_2630; // @[NV_NVDLA_CSC_dl_for_check.scala 1056:29:@1583.4]
  assign _T_2633 = {_T_2444,_T_2444,_T_2444,_T_2444}; // @[Cat.scala 30:58:@1584.4]
  assign _T_2634 = _T_2631 ? 1024'h0 : _T_2633; // @[NV_NVDLA_CSC_dl_for_check.scala 1056:28:@1585.4]
  assign _T_2635 = _T_834[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1586.4]
  assign _T_2636 = ~ _T_2635; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:29:@1587.4]
  assign _T_2639 = _T_2636 ? 1024'h0 : _T_2633; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:28:@1589.4]
  assign _T_2640 = _T_834[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1058:39:@1590.4]
  assign _T_2641 = ~ _T_2640; // @[NV_NVDLA_CSC_dl_for_check.scala 1058:29:@1591.4]
  assign _T_2644 = _T_2641 ? 1024'h0 : _T_2633; // @[NV_NVDLA_CSC_dl_for_check.scala 1058:28:@1593.4]
  assign _T_2646 = {_T_2185,3'h0}; // @[Cat.scala 30:58:@1594.4]
  assign _T_2647 = _T_2629 >> _T_2646; // @[NV_NVDLA_CSC_dl_for_check.scala 1060:41:@1595.4]
  assign _T_2648 = _T_2647[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1060:82:@1596.4]
  assign _T_2650 = {_T_2188,3'h0}; // @[Cat.scala 30:58:@1597.4]
  assign _T_2651 = _T_2634 >> _T_2650; // @[NV_NVDLA_CSC_dl_for_check.scala 1061:41:@1598.4]
  assign _T_2652 = _T_2651[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1061:82:@1599.4]
  assign _T_2654 = {_T_2191,3'h0}; // @[Cat.scala 30:58:@1600.4]
  assign _T_2655 = _T_2639 >> _T_2654; // @[NV_NVDLA_CSC_dl_for_check.scala 1062:41:@1601.4]
  assign _T_2656 = _T_2655[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1062:82:@1602.4]
  assign _T_2658 = {_T_2194,3'h0}; // @[Cat.scala 30:58:@1603.4]
  assign _T_2659 = _T_2644 >> _T_2658; // @[NV_NVDLA_CSC_dl_for_check.scala 1063:41:@1604.4]
  assign _T_2660 = _T_2659[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1063:82:@1605.4]
  assign _T_2661 = _T_834[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:36:@1606.4]
  assign _T_2662 = ~ _T_2661; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:26:@1607.4]
  assign _T_2665 = _T_896 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:41:@1608.4]
  assign _T_2666 = _T_2660[127:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:81:@1609.4]
  assign _T_2672 = {_T_2666,_T_2624,_T_2622,_T_2618}; // @[Cat.scala 30:58:@1615.4]
  assign _T_2674 = _T_896 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1067:41:@1616.4]
  assign _T_2675 = _T_2652[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1067:81:@1617.4]
  assign _T_2677 = {_T_2675,_T_2614}; // @[Cat.scala 30:58:@1619.4]
  assign _T_2679 = _T_2674 ? _T_2677 : _T_2648; // @[NV_NVDLA_CSC_dl_for_check.scala 1067:25:@1621.4]
  assign _T_2680 = _T_2665 ? _T_2672 : _T_2679; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:25:@1622.4]
  assign _T_2681 = _T_2662 ? 512'h0 : _T_2680; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:25:@1623.4]
  assign _T_2752 = _T_2681[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1625.4]
  assign _T_2753 = _T_2681[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1627.4]
  assign _T_2754 = _T_2681[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1629.4]
  assign _T_2755 = _T_2681[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1631.4]
  assign _T_2756 = _T_2681[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1633.4]
  assign _T_2757 = _T_2681[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1635.4]
  assign _T_2758 = _T_2681[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1637.4]
  assign _T_2759 = _T_2681[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1639.4]
  assign _T_2760 = _T_2681[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1641.4]
  assign _T_2761 = _T_2681[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1643.4]
  assign _T_2762 = _T_2681[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1645.4]
  assign _T_2763 = _T_2681[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1647.4]
  assign _T_2764 = _T_2681[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1649.4]
  assign _T_2765 = _T_2681[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1651.4]
  assign _T_2766 = _T_2681[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1653.4]
  assign _T_2767 = _T_2681[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1655.4]
  assign _T_2768 = _T_2681[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1657.4]
  assign _T_2769 = _T_2681[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1659.4]
  assign _T_2770 = _T_2681[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1661.4]
  assign _T_2771 = _T_2681[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1663.4]
  assign _T_2772 = _T_2681[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1665.4]
  assign _T_2773 = _T_2681[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1667.4]
  assign _T_2774 = _T_2681[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1669.4]
  assign _T_2775 = _T_2681[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1671.4]
  assign _T_2776 = _T_2681[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1673.4]
  assign _T_2777 = _T_2681[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1675.4]
  assign _T_2778 = _T_2681[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1677.4]
  assign _T_2779 = _T_2681[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1679.4]
  assign _T_2780 = _T_2681[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1681.4]
  assign _T_2781 = _T_2681[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1683.4]
  assign _T_2782 = _T_2681[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1685.4]
  assign _T_2783 = _T_2681[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1687.4]
  assign _T_2784 = _T_2681[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1689.4]
  assign _T_2785 = _T_2681[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1691.4]
  assign _T_2786 = _T_2681[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1693.4]
  assign _T_2787 = _T_2681[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1695.4]
  assign _T_2788 = _T_2681[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1697.4]
  assign _T_2789 = _T_2681[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1699.4]
  assign _T_2790 = _T_2681[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1701.4]
  assign _T_2791 = _T_2681[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1703.4]
  assign _T_2792 = _T_2681[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1705.4]
  assign _T_2793 = _T_2681[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1707.4]
  assign _T_2794 = _T_2681[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1709.4]
  assign _T_2795 = _T_2681[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1711.4]
  assign _T_2796 = _T_2681[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1713.4]
  assign _T_2797 = _T_2681[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1715.4]
  assign _T_2798 = _T_2681[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1717.4]
  assign _T_2799 = _T_2681[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1719.4]
  assign _T_2800 = _T_2681[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1721.4]
  assign _T_2801 = _T_2681[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1723.4]
  assign _T_2802 = _T_2681[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1725.4]
  assign _T_2803 = _T_2681[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1727.4]
  assign _T_2804 = _T_2681[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1729.4]
  assign _T_2805 = _T_2681[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1731.4]
  assign _T_2806 = _T_2681[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1733.4]
  assign _T_2807 = _T_2681[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1735.4]
  assign _T_2808 = _T_2681[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1737.4]
  assign _T_2809 = _T_2681[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1739.4]
  assign _T_2810 = _T_2681[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1741.4]
  assign _T_2811 = _T_2681[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1743.4]
  assign _T_2812 = _T_2681[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1745.4]
  assign _T_2813 = _T_2681[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1747.4]
  assign _T_2814 = _T_2681[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1749.4]
  assign _T_2815 = _T_2681[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:37:@1751.4]
  assign _T_2817 = _T_899 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:59:@1753.4]
  assign _T_2818 = _T_2211 & _T_2817; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:41:@1754.4]
  assign _T_2820 = _T_899 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:59:@1755.4]
  assign _T_2821 = _T_2214 & _T_2820; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:41:@1756.4]
  assign _T_2824 = _T_2217 & _T_2820; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:41:@1758.4]
  assign _GEN_149 = _T_2818 ? _T_2648 : {{256'd0}, _T_2614}; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:24:@1759.4]
  assign _GEN_150 = _T_2821 ? _T_2614 : {{128'd0}, _T_2616}; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:24:@1762.4]
  assign _GEN_151 = _T_2821 ? _T_2652 : {{384'd0}, _T_2620}; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:24:@1762.4]
  assign _GEN_154 = _T_2824 ? _T_2656 : {{384'd0}, _T_2624}; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:24:@1766.4]
  assign _T_2830 = 319'hffffffffffffffff << _T_2288; // @[NV_NVDLA_CSC_dl_for_check.scala 1096:56:@1772.4]
  assign _T_2831 = _T_2830[63:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1096:73:@1773.4]
  assign _T_2832 = ~ _T_2831; // @[NV_NVDLA_CSC_dl_for_check.scala 1096:24:@1774.4]
  assign _T_2834 = _T_2289 >= 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:51:@1775.4]
  assign _T_2841 = _T_2834 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:32:@1777.4]
  assign _T_2843 = _T_2289 >= 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:51:@1778.4]
  assign _T_2850 = _T_2843 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:32:@1780.4]
  assign _T_2852 = _T_2289 == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:51:@1781.4]
  assign _T_2859 = _T_2852 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:32:@1783.4]
  assign _T_2860 = _T_2841[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:57:@1784.4]
  assign _T_2866 = {_T_2860,32'hffffffff}; // @[Cat.scala 30:58:@1786.4]
  assign _T_2867 = _T_2859[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1103:57:@1787.4]
  assign _T_2868 = _T_2850[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1103:106:@1788.4]
  assign _T_2869 = _T_2841[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1103:155:@1789.4]
  assign _T_2877 = {_T_2867,_T_2868,_T_2869,16'hffff}; // @[Cat.scala 30:58:@1793.4]
  assign _T_2879 = _T_905 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:43:@1794.4]
  assign _T_2880 = _T_2832[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:89:@1795.4]
  assign _T_2882 = {_T_2880,_T_2880,_T_2880,_T_2880}; // @[Cat.scala 30:58:@1797.4]
  assign _T_2883 = _T_2882 & _T_2877; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:116:@1798.4]
  assign _T_2885 = _T_905 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:43:@1799.4]
  assign _T_2886 = _T_2832[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:89:@1800.4]
  assign _T_2887 = {_T_2886,_T_2886}; // @[Cat.scala 30:58:@1801.4]
  assign _T_2888 = _T_2887 & _T_2866; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:116:@1802.4]
  assign _T_2889 = _T_2885 ? _T_2888 : _T_2832; // @[NV_NVDLA_CSC_dl_for_check.scala 1106:26:@1803.4]
  assign _T_2890 = _T_2879 ? _T_2883 : _T_2889; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:26:@1804.4]
  assign _T_2891 = _T_834[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:35:@1805.4]
  assign _T_2892_0 = _T_2891 ? _T_2752 : _T_2549; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_1 = _T_2891 ? _T_2753 : _T_2550; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_2 = _T_2891 ? _T_2754 : _T_2551; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_3 = _T_2891 ? _T_2755 : _T_2552; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_4 = _T_2891 ? _T_2756 : _T_2553; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_5 = _T_2891 ? _T_2757 : _T_2554; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_6 = _T_2891 ? _T_2758 : _T_2555; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_7 = _T_2891 ? _T_2759 : _T_2556; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_8 = _T_2891 ? _T_2760 : _T_2557; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_9 = _T_2891 ? _T_2761 : _T_2558; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_10 = _T_2891 ? _T_2762 : _T_2559; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_11 = _T_2891 ? _T_2763 : _T_2560; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_12 = _T_2891 ? _T_2764 : _T_2561; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_13 = _T_2891 ? _T_2765 : _T_2562; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_14 = _T_2891 ? _T_2766 : _T_2563; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_15 = _T_2891 ? _T_2767 : _T_2564; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_16 = _T_2891 ? _T_2768 : _T_2565; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_17 = _T_2891 ? _T_2769 : _T_2566; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_18 = _T_2891 ? _T_2770 : _T_2567; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_19 = _T_2891 ? _T_2771 : _T_2568; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_20 = _T_2891 ? _T_2772 : _T_2569; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_21 = _T_2891 ? _T_2773 : _T_2570; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_22 = _T_2891 ? _T_2774 : _T_2571; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_23 = _T_2891 ? _T_2775 : _T_2572; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_24 = _T_2891 ? _T_2776 : _T_2573; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_25 = _T_2891 ? _T_2777 : _T_2574; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_26 = _T_2891 ? _T_2778 : _T_2575; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_27 = _T_2891 ? _T_2779 : _T_2576; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_28 = _T_2891 ? _T_2780 : _T_2577; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_29 = _T_2891 ? _T_2781 : _T_2578; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_30 = _T_2891 ? _T_2782 : _T_2579; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_31 = _T_2891 ? _T_2783 : _T_2580; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_32 = _T_2891 ? _T_2784 : _T_2581; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_33 = _T_2891 ? _T_2785 : _T_2582; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_34 = _T_2891 ? _T_2786 : _T_2583; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_35 = _T_2891 ? _T_2787 : _T_2584; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_36 = _T_2891 ? _T_2788 : _T_2585; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_37 = _T_2891 ? _T_2789 : _T_2586; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_38 = _T_2891 ? _T_2790 : _T_2587; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_39 = _T_2891 ? _T_2791 : _T_2588; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_40 = _T_2891 ? _T_2792 : _T_2589; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_41 = _T_2891 ? _T_2793 : _T_2590; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_42 = _T_2891 ? _T_2794 : _T_2591; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_43 = _T_2891 ? _T_2795 : _T_2592; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_44 = _T_2891 ? _T_2796 : _T_2593; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_45 = _T_2891 ? _T_2797 : _T_2594; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_46 = _T_2891 ? _T_2798 : _T_2595; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_47 = _T_2891 ? _T_2799 : _T_2596; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_48 = _T_2891 ? _T_2800 : _T_2597; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_49 = _T_2891 ? _T_2801 : _T_2598; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_50 = _T_2891 ? _T_2802 : _T_2599; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_51 = _T_2891 ? _T_2803 : _T_2600; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_52 = _T_2891 ? _T_2804 : _T_2601; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_53 = _T_2891 ? _T_2805 : _T_2602; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_54 = _T_2891 ? _T_2806 : _T_2603; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_55 = _T_2891 ? _T_2807 : _T_2604; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_56 = _T_2891 ? _T_2808 : _T_2605; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_57 = _T_2891 ? _T_2809 : _T_2606; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_58 = _T_2891 ? _T_2810 : _T_2607; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_59 = _T_2891 ? _T_2811 : _T_2608; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_60 = _T_2891 ? _T_2812 : _T_2609; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_61 = _T_2891 ? _T_2813 : _T_2610; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_62 = _T_2891 ? _T_2814 : _T_2611; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_2892_63 = _T_2891 ? _T_2815 : _T_2612; // @[NV_NVDLA_CSC_dl_for_check.scala 1110:25:@1806.4]
  assign _T_3025 = _T_2892_0 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1807.4]
  assign _T_3027 = _T_2892_1 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1808.4]
  assign _T_3029 = _T_2892_2 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1809.4]
  assign _T_3031 = _T_2892_3 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1810.4]
  assign _T_3033 = _T_2892_4 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1811.4]
  assign _T_3035 = _T_2892_5 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1812.4]
  assign _T_3037 = _T_2892_6 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1813.4]
  assign _T_3039 = _T_2892_7 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1814.4]
  assign _T_3041 = _T_2892_8 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1815.4]
  assign _T_3043 = _T_2892_9 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1816.4]
  assign _T_3045 = _T_2892_10 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1817.4]
  assign _T_3047 = _T_2892_11 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1818.4]
  assign _T_3049 = _T_2892_12 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1819.4]
  assign _T_3051 = _T_2892_13 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1820.4]
  assign _T_3053 = _T_2892_14 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1821.4]
  assign _T_3055 = _T_2892_15 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1822.4]
  assign _T_3057 = _T_2892_16 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1823.4]
  assign _T_3059 = _T_2892_17 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1824.4]
  assign _T_3061 = _T_2892_18 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1825.4]
  assign _T_3063 = _T_2892_19 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1826.4]
  assign _T_3065 = _T_2892_20 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1827.4]
  assign _T_3067 = _T_2892_21 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1828.4]
  assign _T_3069 = _T_2892_22 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1829.4]
  assign _T_3071 = _T_2892_23 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1830.4]
  assign _T_3073 = _T_2892_24 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1831.4]
  assign _T_3075 = _T_2892_25 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1832.4]
  assign _T_3077 = _T_2892_26 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1833.4]
  assign _T_3079 = _T_2892_27 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1834.4]
  assign _T_3081 = _T_2892_28 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1835.4]
  assign _T_3083 = _T_2892_29 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1836.4]
  assign _T_3085 = _T_2892_30 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1837.4]
  assign _T_3087 = _T_2892_31 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1838.4]
  assign _T_3089 = _T_2892_32 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1839.4]
  assign _T_3091 = _T_2892_33 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1840.4]
  assign _T_3093 = _T_2892_34 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1841.4]
  assign _T_3095 = _T_2892_35 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1842.4]
  assign _T_3097 = _T_2892_36 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1843.4]
  assign _T_3099 = _T_2892_37 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1844.4]
  assign _T_3101 = _T_2892_38 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1845.4]
  assign _T_3103 = _T_2892_39 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1846.4]
  assign _T_3105 = _T_2892_40 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1847.4]
  assign _T_3107 = _T_2892_41 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1848.4]
  assign _T_3109 = _T_2892_42 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1849.4]
  assign _T_3111 = _T_2892_43 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1850.4]
  assign _T_3113 = _T_2892_44 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1851.4]
  assign _T_3115 = _T_2892_45 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1852.4]
  assign _T_3117 = _T_2892_46 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1853.4]
  assign _T_3119 = _T_2892_47 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1854.4]
  assign _T_3121 = _T_2892_48 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1855.4]
  assign _T_3123 = _T_2892_49 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1856.4]
  assign _T_3125 = _T_2892_50 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1857.4]
  assign _T_3127 = _T_2892_51 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1858.4]
  assign _T_3129 = _T_2892_52 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1859.4]
  assign _T_3131 = _T_2892_53 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1860.4]
  assign _T_3133 = _T_2892_54 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1861.4]
  assign _T_3135 = _T_2892_55 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1862.4]
  assign _T_3137 = _T_2892_56 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1863.4]
  assign _T_3139 = _T_2892_57 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1864.4]
  assign _T_3141 = _T_2892_58 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1865.4]
  assign _T_3143 = _T_2892_59 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1866.4]
  assign _T_3145 = _T_2892_60 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1867.4]
  assign _T_3147 = _T_2892_61 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1868.4]
  assign _T_3149 = _T_2892_62 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1869.4]
  assign _T_3151 = _T_2892_63 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:97:@1870.4]
  assign _T_3222 = _T_2890[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1936.4]
  assign _T_3223 = _T_3222 & _T_3025; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1937.4]
  assign _T_3224 = _T_2890[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1938.4]
  assign _T_3225 = _T_3224 & _T_3027; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1939.4]
  assign _T_3226 = _T_2890[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1940.4]
  assign _T_3227 = _T_3226 & _T_3029; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1941.4]
  assign _T_3228 = _T_2890[3]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1942.4]
  assign _T_3229 = _T_3228 & _T_3031; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1943.4]
  assign _T_3230 = _T_2890[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1944.4]
  assign _T_3231 = _T_3230 & _T_3033; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1945.4]
  assign _T_3232 = _T_2890[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1946.4]
  assign _T_3233 = _T_3232 & _T_3035; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1947.4]
  assign _T_3234 = _T_2890[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1948.4]
  assign _T_3235 = _T_3234 & _T_3037; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1949.4]
  assign _T_3236 = _T_2890[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1950.4]
  assign _T_3237 = _T_3236 & _T_3039; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1951.4]
  assign _T_3238 = _T_2890[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1952.4]
  assign _T_3239 = _T_3238 & _T_3041; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1953.4]
  assign _T_3240 = _T_2890[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1954.4]
  assign _T_3241 = _T_3240 & _T_3043; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1955.4]
  assign _T_3242 = _T_2890[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1956.4]
  assign _T_3243 = _T_3242 & _T_3045; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1957.4]
  assign _T_3244 = _T_2890[11]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1958.4]
  assign _T_3245 = _T_3244 & _T_3047; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1959.4]
  assign _T_3246 = _T_2890[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1960.4]
  assign _T_3247 = _T_3246 & _T_3049; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1961.4]
  assign _T_3248 = _T_2890[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1962.4]
  assign _T_3249 = _T_3248 & _T_3051; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1963.4]
  assign _T_3250 = _T_2890[14]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1964.4]
  assign _T_3251 = _T_3250 & _T_3053; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1965.4]
  assign _T_3252 = _T_2890[15]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1966.4]
  assign _T_3253 = _T_3252 & _T_3055; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1967.4]
  assign _T_3254 = _T_2890[16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1968.4]
  assign _T_3255 = _T_3254 & _T_3057; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1969.4]
  assign _T_3256 = _T_2890[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1970.4]
  assign _T_3257 = _T_3256 & _T_3059; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1971.4]
  assign _T_3258 = _T_2890[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1972.4]
  assign _T_3259 = _T_3258 & _T_3061; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1973.4]
  assign _T_3260 = _T_2890[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1974.4]
  assign _T_3261 = _T_3260 & _T_3063; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1975.4]
  assign _T_3262 = _T_2890[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1976.4]
  assign _T_3263 = _T_3262 & _T_3065; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1977.4]
  assign _T_3264 = _T_2890[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1978.4]
  assign _T_3265 = _T_3264 & _T_3067; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1979.4]
  assign _T_3266 = _T_2890[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1980.4]
  assign _T_3267 = _T_3266 & _T_3069; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1981.4]
  assign _T_3268 = _T_2890[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1982.4]
  assign _T_3269 = _T_3268 & _T_3071; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1983.4]
  assign _T_3270 = _T_2890[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1984.4]
  assign _T_3271 = _T_3270 & _T_3073; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1985.4]
  assign _T_3272 = _T_2890[25]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1986.4]
  assign _T_3273 = _T_3272 & _T_3075; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1987.4]
  assign _T_3274 = _T_2890[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1988.4]
  assign _T_3275 = _T_3274 & _T_3077; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1989.4]
  assign _T_3276 = _T_2890[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1990.4]
  assign _T_3277 = _T_3276 & _T_3079; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1991.4]
  assign _T_3278 = _T_2890[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1992.4]
  assign _T_3279 = _T_3278 & _T_3081; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1993.4]
  assign _T_3280 = _T_2890[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1994.4]
  assign _T_3281 = _T_3280 & _T_3083; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1995.4]
  assign _T_3282 = _T_2890[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1996.4]
  assign _T_3283 = _T_3282 & _T_3085; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1997.4]
  assign _T_3284 = _T_2890[31]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@1998.4]
  assign _T_3285 = _T_3284 & _T_3087; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@1999.4]
  assign _T_3286 = _T_2890[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2000.4]
  assign _T_3287 = _T_3286 & _T_3089; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2001.4]
  assign _T_3288 = _T_2890[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2002.4]
  assign _T_3289 = _T_3288 & _T_3091; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2003.4]
  assign _T_3290 = _T_2890[34]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2004.4]
  assign _T_3291 = _T_3290 & _T_3093; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2005.4]
  assign _T_3292 = _T_2890[35]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2006.4]
  assign _T_3293 = _T_3292 & _T_3095; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2007.4]
  assign _T_3294 = _T_2890[36]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2008.4]
  assign _T_3295 = _T_3294 & _T_3097; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2009.4]
  assign _T_3296 = _T_2890[37]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2010.4]
  assign _T_3297 = _T_3296 & _T_3099; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2011.4]
  assign _T_3298 = _T_2890[38]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2012.4]
  assign _T_3299 = _T_3298 & _T_3101; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2013.4]
  assign _T_3300 = _T_2890[39]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2014.4]
  assign _T_3301 = _T_3300 & _T_3103; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2015.4]
  assign _T_3302 = _T_2890[40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2016.4]
  assign _T_3303 = _T_3302 & _T_3105; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2017.4]
  assign _T_3304 = _T_2890[41]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2018.4]
  assign _T_3305 = _T_3304 & _T_3107; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2019.4]
  assign _T_3306 = _T_2890[42]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2020.4]
  assign _T_3307 = _T_3306 & _T_3109; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2021.4]
  assign _T_3308 = _T_2890[43]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2022.4]
  assign _T_3309 = _T_3308 & _T_3111; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2023.4]
  assign _T_3310 = _T_2890[44]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2024.4]
  assign _T_3311 = _T_3310 & _T_3113; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2025.4]
  assign _T_3312 = _T_2890[45]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2026.4]
  assign _T_3313 = _T_3312 & _T_3115; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2027.4]
  assign _T_3314 = _T_2890[46]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2028.4]
  assign _T_3315 = _T_3314 & _T_3117; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2029.4]
  assign _T_3316 = _T_2890[47]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2030.4]
  assign _T_3317 = _T_3316 & _T_3119; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2031.4]
  assign _T_3318 = _T_2890[48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2032.4]
  assign _T_3319 = _T_3318 & _T_3121; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2033.4]
  assign _T_3320 = _T_2890[49]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2034.4]
  assign _T_3321 = _T_3320 & _T_3123; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2035.4]
  assign _T_3322 = _T_2890[50]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2036.4]
  assign _T_3323 = _T_3322 & _T_3125; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2037.4]
  assign _T_3324 = _T_2890[51]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2038.4]
  assign _T_3325 = _T_3324 & _T_3127; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2039.4]
  assign _T_3326 = _T_2890[52]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2040.4]
  assign _T_3327 = _T_3326 & _T_3129; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2041.4]
  assign _T_3328 = _T_2890[53]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2042.4]
  assign _T_3329 = _T_3328 & _T_3131; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2043.4]
  assign _T_3330 = _T_2890[54]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2044.4]
  assign _T_3331 = _T_3330 & _T_3133; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2045.4]
  assign _T_3332 = _T_2890[55]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2046.4]
  assign _T_3333 = _T_3332 & _T_3135; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2047.4]
  assign _T_3334 = _T_2890[56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2048.4]
  assign _T_3335 = _T_3334 & _T_3137; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2049.4]
  assign _T_3336 = _T_2890[57]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2050.4]
  assign _T_3337 = _T_3336 & _T_3139; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2051.4]
  assign _T_3338 = _T_2890[58]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2052.4]
  assign _T_3339 = _T_3338 & _T_3141; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2053.4]
  assign _T_3340 = _T_2890[59]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2054.4]
  assign _T_3341 = _T_3340 & _T_3143; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2055.4]
  assign _T_3342 = _T_2890[60]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2056.4]
  assign _T_3343 = _T_3342 & _T_3145; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2057.4]
  assign _T_3344 = _T_2890[61]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2058.4]
  assign _T_3345 = _T_3344 & _T_3147; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2059.4]
  assign _T_3346 = _T_2890[62]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2060.4]
  assign _T_3347 = _T_3346 & _T_3149; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2061.4]
  assign _T_3348 = _T_2890[63]; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:80:@2062.4]
  assign _T_3349 = _T_3348 & _T_3151; // @[NV_NVDLA_CSC_dl_for_check.scala 1112:83:@2063.4]
  assign _GEN_156 = _T_2251 ? _T_3223 : _T_3692_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_157 = _T_2251 ? _T_3225 : _T_3692_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_158 = _T_2251 ? _T_3227 : _T_3692_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_159 = _T_2251 ? _T_3229 : _T_3692_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_160 = _T_2251 ? _T_3231 : _T_3692_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_161 = _T_2251 ? _T_3233 : _T_3692_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_162 = _T_2251 ? _T_3235 : _T_3692_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_163 = _T_2251 ? _T_3237 : _T_3692_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_164 = _T_2251 ? _T_3239 : _T_3692_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_165 = _T_2251 ? _T_3241 : _T_3692_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_166 = _T_2251 ? _T_3243 : _T_3692_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_167 = _T_2251 ? _T_3245 : _T_3692_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_168 = _T_2251 ? _T_3247 : _T_3692_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_169 = _T_2251 ? _T_3249 : _T_3692_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_170 = _T_2251 ? _T_3251 : _T_3692_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_171 = _T_2251 ? _T_3253 : _T_3692_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_172 = _T_2251 ? _T_3255 : _T_3692_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_173 = _T_2251 ? _T_3257 : _T_3692_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_174 = _T_2251 ? _T_3259 : _T_3692_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_175 = _T_2251 ? _T_3261 : _T_3692_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_176 = _T_2251 ? _T_3263 : _T_3692_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_177 = _T_2251 ? _T_3265 : _T_3692_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_178 = _T_2251 ? _T_3267 : _T_3692_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_179 = _T_2251 ? _T_3269 : _T_3692_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_180 = _T_2251 ? _T_3271 : _T_3692_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_181 = _T_2251 ? _T_3273 : _T_3692_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_182 = _T_2251 ? _T_3275 : _T_3692_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_183 = _T_2251 ? _T_3277 : _T_3692_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_184 = _T_2251 ? _T_3279 : _T_3692_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_185 = _T_2251 ? _T_3281 : _T_3692_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_186 = _T_2251 ? _T_3283 : _T_3692_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_187 = _T_2251 ? _T_3285 : _T_3692_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_188 = _T_2251 ? _T_3287 : _T_3692_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_189 = _T_2251 ? _T_3289 : _T_3692_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_190 = _T_2251 ? _T_3291 : _T_3692_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_191 = _T_2251 ? _T_3293 : _T_3692_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_192 = _T_2251 ? _T_3295 : _T_3692_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_193 = _T_2251 ? _T_3297 : _T_3692_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_194 = _T_2251 ? _T_3299 : _T_3692_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_195 = _T_2251 ? _T_3301 : _T_3692_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_196 = _T_2251 ? _T_3303 : _T_3692_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_197 = _T_2251 ? _T_3305 : _T_3692_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_198 = _T_2251 ? _T_3307 : _T_3692_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_199 = _T_2251 ? _T_3309 : _T_3692_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_200 = _T_2251 ? _T_3311 : _T_3692_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_201 = _T_2251 ? _T_3313 : _T_3692_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_202 = _T_2251 ? _T_3315 : _T_3692_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_203 = _T_2251 ? _T_3317 : _T_3692_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_204 = _T_2251 ? _T_3319 : _T_3692_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_205 = _T_2251 ? _T_3321 : _T_3692_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_206 = _T_2251 ? _T_3323 : _T_3692_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_207 = _T_2251 ? _T_3325 : _T_3692_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_208 = _T_2251 ? _T_3327 : _T_3692_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_209 = _T_2251 ? _T_3329 : _T_3692_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_210 = _T_2251 ? _T_3331 : _T_3692_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_211 = _T_2251 ? _T_3333 : _T_3692_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_212 = _T_2251 ? _T_3335 : _T_3692_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_213 = _T_2251 ? _T_3337 : _T_3692_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_214 = _T_2251 ? _T_3339 : _T_3692_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_215 = _T_2251 ? _T_3341 : _T_3692_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_216 = _T_2251 ? _T_3343 : _T_3692_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_217 = _T_2251 ? _T_3345 : _T_3692_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_218 = _T_2251 ? _T_3347 : _T_3692_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _GEN_219 = _T_2251 ? _T_3349 : _T_3692_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:30:@2202.4]
  assign _T_3959 = _T_2251 & _T_3223; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2268.4]
  assign _T_3960 = _T_2251 & _T_3225; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2272.4]
  assign _T_3961 = _T_2251 & _T_3227; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2276.4]
  assign _T_3962 = _T_2251 & _T_3229; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2280.4]
  assign _T_3963 = _T_2251 & _T_3231; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2284.4]
  assign _T_3964 = _T_2251 & _T_3233; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2288.4]
  assign _T_3965 = _T_2251 & _T_3235; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2292.4]
  assign _T_3966 = _T_2251 & _T_3237; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2296.4]
  assign _T_3967 = _T_2251 & _T_3239; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2300.4]
  assign _T_3968 = _T_2251 & _T_3241; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2304.4]
  assign _T_3969 = _T_2251 & _T_3243; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2308.4]
  assign _T_3970 = _T_2251 & _T_3245; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2312.4]
  assign _T_3971 = _T_2251 & _T_3247; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2316.4]
  assign _T_3972 = _T_2251 & _T_3249; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2320.4]
  assign _T_3973 = _T_2251 & _T_3251; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2324.4]
  assign _T_3974 = _T_2251 & _T_3253; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2328.4]
  assign _T_3975 = _T_2251 & _T_3255; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2332.4]
  assign _T_3976 = _T_2251 & _T_3257; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2336.4]
  assign _T_3977 = _T_2251 & _T_3259; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2340.4]
  assign _T_3978 = _T_2251 & _T_3261; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2344.4]
  assign _T_3979 = _T_2251 & _T_3263; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2348.4]
  assign _T_3980 = _T_2251 & _T_3265; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2352.4]
  assign _T_3981 = _T_2251 & _T_3267; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2356.4]
  assign _T_3982 = _T_2251 & _T_3269; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2360.4]
  assign _T_3983 = _T_2251 & _T_3271; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2364.4]
  assign _T_3984 = _T_2251 & _T_3273; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2368.4]
  assign _T_3985 = _T_2251 & _T_3275; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2372.4]
  assign _T_3986 = _T_2251 & _T_3277; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2376.4]
  assign _T_3987 = _T_2251 & _T_3279; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2380.4]
  assign _T_3988 = _T_2251 & _T_3281; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2384.4]
  assign _T_3989 = _T_2251 & _T_3283; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2388.4]
  assign _T_3990 = _T_2251 & _T_3285; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2392.4]
  assign _T_3991 = _T_2251 & _T_3287; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2396.4]
  assign _T_3992 = _T_2251 & _T_3289; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2400.4]
  assign _T_3993 = _T_2251 & _T_3291; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2404.4]
  assign _T_3994 = _T_2251 & _T_3293; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2408.4]
  assign _T_3995 = _T_2251 & _T_3295; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2412.4]
  assign _T_3996 = _T_2251 & _T_3297; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2416.4]
  assign _T_3997 = _T_2251 & _T_3299; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2420.4]
  assign _T_3998 = _T_2251 & _T_3301; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2424.4]
  assign _T_3999 = _T_2251 & _T_3303; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2428.4]
  assign _T_4000 = _T_2251 & _T_3305; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2432.4]
  assign _T_4001 = _T_2251 & _T_3307; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2436.4]
  assign _T_4002 = _T_2251 & _T_3309; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2440.4]
  assign _T_4003 = _T_2251 & _T_3311; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2444.4]
  assign _T_4004 = _T_2251 & _T_3313; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2448.4]
  assign _T_4005 = _T_2251 & _T_3315; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2452.4]
  assign _T_4006 = _T_2251 & _T_3317; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2456.4]
  assign _T_4007 = _T_2251 & _T_3319; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2460.4]
  assign _T_4008 = _T_2251 & _T_3321; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2464.4]
  assign _T_4009 = _T_2251 & _T_3323; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2468.4]
  assign _T_4010 = _T_2251 & _T_3325; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2472.4]
  assign _T_4011 = _T_2251 & _T_3327; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2476.4]
  assign _T_4012 = _T_2251 & _T_3329; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2480.4]
  assign _T_4013 = _T_2251 & _T_3331; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2484.4]
  assign _T_4014 = _T_2251 & _T_3333; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2488.4]
  assign _T_4015 = _T_2251 & _T_3335; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2492.4]
  assign _T_4016 = _T_2251 & _T_3337; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2496.4]
  assign _T_4017 = _T_2251 & _T_3339; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2500.4]
  assign _T_4018 = _T_2251 & _T_3341; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2504.4]
  assign _T_4019 = _T_2251 & _T_3343; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2508.4]
  assign _T_4020 = _T_2251 & _T_3345; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2512.4]
  assign _T_4021 = _T_2251 & _T_3347; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2516.4]
  assign _T_4022 = _T_2251 & _T_3349; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:34:@2520.4]
  assign _T_4562 = ~ _T_3422; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:24:@2593.4]
  assign _T_4697_0 = _T_4562 ? 1'h0 : _T_3692_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_1 = _T_4562 ? 1'h0 : _T_3692_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_2 = _T_4562 ? 1'h0 : _T_3692_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_3 = _T_4562 ? 1'h0 : _T_3692_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_4 = _T_4562 ? 1'h0 : _T_3692_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_5 = _T_4562 ? 1'h0 : _T_3692_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_6 = _T_4562 ? 1'h0 : _T_3692_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_7 = _T_4562 ? 1'h0 : _T_3692_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_8 = _T_4562 ? 1'h0 : _T_3692_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_9 = _T_4562 ? 1'h0 : _T_3692_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_10 = _T_4562 ? 1'h0 : _T_3692_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_11 = _T_4562 ? 1'h0 : _T_3692_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_12 = _T_4562 ? 1'h0 : _T_3692_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_13 = _T_4562 ? 1'h0 : _T_3692_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_14 = _T_4562 ? 1'h0 : _T_3692_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_15 = _T_4562 ? 1'h0 : _T_3692_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_16 = _T_4562 ? 1'h0 : _T_3692_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_17 = _T_4562 ? 1'h0 : _T_3692_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_18 = _T_4562 ? 1'h0 : _T_3692_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_19 = _T_4562 ? 1'h0 : _T_3692_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_20 = _T_4562 ? 1'h0 : _T_3692_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_21 = _T_4562 ? 1'h0 : _T_3692_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_22 = _T_4562 ? 1'h0 : _T_3692_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_23 = _T_4562 ? 1'h0 : _T_3692_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_24 = _T_4562 ? 1'h0 : _T_3692_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_25 = _T_4562 ? 1'h0 : _T_3692_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_26 = _T_4562 ? 1'h0 : _T_3692_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_27 = _T_4562 ? 1'h0 : _T_3692_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_28 = _T_4562 ? 1'h0 : _T_3692_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_29 = _T_4562 ? 1'h0 : _T_3692_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_30 = _T_4562 ? 1'h0 : _T_3692_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_31 = _T_4562 ? 1'h0 : _T_3692_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_32 = _T_4562 ? 1'h0 : _T_3692_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_33 = _T_4562 ? 1'h0 : _T_3692_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_34 = _T_4562 ? 1'h0 : _T_3692_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_35 = _T_4562 ? 1'h0 : _T_3692_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_36 = _T_4562 ? 1'h0 : _T_3692_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_37 = _T_4562 ? 1'h0 : _T_3692_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_38 = _T_4562 ? 1'h0 : _T_3692_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_39 = _T_4562 ? 1'h0 : _T_3692_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_40 = _T_4562 ? 1'h0 : _T_3692_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_41 = _T_4562 ? 1'h0 : _T_3692_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_42 = _T_4562 ? 1'h0 : _T_3692_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_43 = _T_4562 ? 1'h0 : _T_3692_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_44 = _T_4562 ? 1'h0 : _T_3692_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_45 = _T_4562 ? 1'h0 : _T_3692_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_46 = _T_4562 ? 1'h0 : _T_3692_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_47 = _T_4562 ? 1'h0 : _T_3692_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_48 = _T_4562 ? 1'h0 : _T_3692_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_49 = _T_4562 ? 1'h0 : _T_3692_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_50 = _T_4562 ? 1'h0 : _T_3692_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_51 = _T_4562 ? 1'h0 : _T_3692_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_52 = _T_4562 ? 1'h0 : _T_3692_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_53 = _T_4562 ? 1'h0 : _T_3692_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_54 = _T_4562 ? 1'h0 : _T_3692_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_55 = _T_4562 ? 1'h0 : _T_3692_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_56 = _T_4562 ? 1'h0 : _T_3692_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_57 = _T_4562 ? 1'h0 : _T_3692_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_58 = _T_4562 ? 1'h0 : _T_3692_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_59 = _T_4562 ? 1'h0 : _T_3692_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_60 = _T_4562 ? 1'h0 : _T_3692_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_61 = _T_4562 ? 1'h0 : _T_3692_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_62 = _T_4562 ? 1'h0 : _T_3692_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4697_63 = _T_4562 ? 1'h0 : _T_3692_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:23:@2659.4]
  assign _T_4829 = _T_3422 | _T_4025; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:19:@2661.4]
  assign _GEN_284 = _T_4829 ? _T_4697_0 : _T_4292_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_285 = _T_4829 ? _T_4697_1 : _T_4292_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_286 = _T_4829 ? _T_4697_2 : _T_4292_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_287 = _T_4829 ? _T_4697_3 : _T_4292_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_288 = _T_4829 ? _T_4697_4 : _T_4292_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_289 = _T_4829 ? _T_4697_5 : _T_4292_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_290 = _T_4829 ? _T_4697_6 : _T_4292_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_291 = _T_4829 ? _T_4697_7 : _T_4292_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_292 = _T_4829 ? _T_4697_8 : _T_4292_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_293 = _T_4829 ? _T_4697_9 : _T_4292_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_294 = _T_4829 ? _T_4697_10 : _T_4292_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_295 = _T_4829 ? _T_4697_11 : _T_4292_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_296 = _T_4829 ? _T_4697_12 : _T_4292_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_297 = _T_4829 ? _T_4697_13 : _T_4292_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_298 = _T_4829 ? _T_4697_14 : _T_4292_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_299 = _T_4829 ? _T_4697_15 : _T_4292_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_300 = _T_4829 ? _T_4697_16 : _T_4292_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_301 = _T_4829 ? _T_4697_17 : _T_4292_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_302 = _T_4829 ? _T_4697_18 : _T_4292_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_303 = _T_4829 ? _T_4697_19 : _T_4292_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_304 = _T_4829 ? _T_4697_20 : _T_4292_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_305 = _T_4829 ? _T_4697_21 : _T_4292_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_306 = _T_4829 ? _T_4697_22 : _T_4292_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_307 = _T_4829 ? _T_4697_23 : _T_4292_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_308 = _T_4829 ? _T_4697_24 : _T_4292_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_309 = _T_4829 ? _T_4697_25 : _T_4292_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_310 = _T_4829 ? _T_4697_26 : _T_4292_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_311 = _T_4829 ? _T_4697_27 : _T_4292_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_312 = _T_4829 ? _T_4697_28 : _T_4292_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_313 = _T_4829 ? _T_4697_29 : _T_4292_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_314 = _T_4829 ? _T_4697_30 : _T_4292_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_315 = _T_4829 ? _T_4697_31 : _T_4292_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_316 = _T_4829 ? _T_4697_32 : _T_4292_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_317 = _T_4829 ? _T_4697_33 : _T_4292_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_318 = _T_4829 ? _T_4697_34 : _T_4292_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_319 = _T_4829 ? _T_4697_35 : _T_4292_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_320 = _T_4829 ? _T_4697_36 : _T_4292_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_321 = _T_4829 ? _T_4697_37 : _T_4292_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_322 = _T_4829 ? _T_4697_38 : _T_4292_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_323 = _T_4829 ? _T_4697_39 : _T_4292_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_324 = _T_4829 ? _T_4697_40 : _T_4292_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_325 = _T_4829 ? _T_4697_41 : _T_4292_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_326 = _T_4829 ? _T_4697_42 : _T_4292_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_327 = _T_4829 ? _T_4697_43 : _T_4292_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_328 = _T_4829 ? _T_4697_44 : _T_4292_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_329 = _T_4829 ? _T_4697_45 : _T_4292_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_330 = _T_4829 ? _T_4697_46 : _T_4292_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_331 = _T_4829 ? _T_4697_47 : _T_4292_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_332 = _T_4829 ? _T_4697_48 : _T_4292_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_333 = _T_4829 ? _T_4697_49 : _T_4292_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_334 = _T_4829 ? _T_4697_50 : _T_4292_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_335 = _T_4829 ? _T_4697_51 : _T_4292_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_336 = _T_4829 ? _T_4697_52 : _T_4292_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_337 = _T_4829 ? _T_4697_53 : _T_4292_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_338 = _T_4829 ? _T_4697_54 : _T_4292_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_339 = _T_4829 ? _T_4697_55 : _T_4292_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_340 = _T_4829 ? _T_4697_56 : _T_4292_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_341 = _T_4829 ? _T_4697_57 : _T_4292_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_342 = _T_4829 ? _T_4697_58 : _T_4292_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_343 = _T_4829 ? _T_4697_59 : _T_4292_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_344 = _T_4829 ? _T_4697_60 : _T_4292_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_345 = _T_4829 ? _T_4697_61 : _T_4292_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_346 = _T_4829 ? _T_4697_62 : _T_4292_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_347 = _T_4829 ? _T_4697_63 : _T_4292_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:33:@2662.4]
  assign _GEN_348 = _T_3422 ? {{8'd0}, _T_3422} : _T_4491; // @[NV_NVDLA_CSC_dl_for_check.scala 1160:19:@2728.4]
  assign _T_4833 = ~ _T_4025; // @[NV_NVDLA_CSC_dl_for_check.scala 1174:27:@2925.4]
  assign _T_4835 = _T_4833 ? 9'h0 : _T_4491; // @[NV_NVDLA_CSC_dl_for_check.scala 1174:26:@2926.4]
  assign _T_4843 = _T_4025 | _T_4832; // @[NV_NVDLA_CSC_dl_for_check.scala 1178:85:@2933.4]
  assign _GEN_413 = _T_4843 ? _T_4835 : _T_4845; // @[Reg.scala 20:19:@2935.4]
  assign _GEN_414 = _T_4843 ? _T_4835 : _T_4849; // @[Reg.scala 20:19:@2941.4]
  assign _GEN_415 = _T_4843 ? _T_4292_0 : _T_5117_0; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_416 = _T_4843 ? _T_4292_1 : _T_5117_1; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_417 = _T_4843 ? _T_4292_2 : _T_5117_2; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_418 = _T_4843 ? _T_4292_3 : _T_5117_3; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_419 = _T_4843 ? _T_4292_4 : _T_5117_4; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_420 = _T_4843 ? _T_4292_5 : _T_5117_5; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_421 = _T_4843 ? _T_4292_6 : _T_5117_6; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_422 = _T_4843 ? _T_4292_7 : _T_5117_7; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_423 = _T_4843 ? _T_4292_8 : _T_5117_8; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_424 = _T_4843 ? _T_4292_9 : _T_5117_9; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_425 = _T_4843 ? _T_4292_10 : _T_5117_10; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_426 = _T_4843 ? _T_4292_11 : _T_5117_11; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_427 = _T_4843 ? _T_4292_12 : _T_5117_12; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_428 = _T_4843 ? _T_4292_13 : _T_5117_13; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_429 = _T_4843 ? _T_4292_14 : _T_5117_14; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_430 = _T_4843 ? _T_4292_15 : _T_5117_15; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_431 = _T_4843 ? _T_4292_16 : _T_5117_16; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_432 = _T_4843 ? _T_4292_17 : _T_5117_17; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_433 = _T_4843 ? _T_4292_18 : _T_5117_18; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_434 = _T_4843 ? _T_4292_19 : _T_5117_19; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_435 = _T_4843 ? _T_4292_20 : _T_5117_20; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_436 = _T_4843 ? _T_4292_21 : _T_5117_21; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_437 = _T_4843 ? _T_4292_22 : _T_5117_22; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_438 = _T_4843 ? _T_4292_23 : _T_5117_23; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_439 = _T_4843 ? _T_4292_24 : _T_5117_24; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_440 = _T_4843 ? _T_4292_25 : _T_5117_25; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_441 = _T_4843 ? _T_4292_26 : _T_5117_26; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_442 = _T_4843 ? _T_4292_27 : _T_5117_27; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_443 = _T_4843 ? _T_4292_28 : _T_5117_28; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_444 = _T_4843 ? _T_4292_29 : _T_5117_29; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_445 = _T_4843 ? _T_4292_30 : _T_5117_30; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_446 = _T_4843 ? _T_4292_31 : _T_5117_31; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_447 = _T_4843 ? _T_4292_32 : _T_5117_32; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_448 = _T_4843 ? _T_4292_33 : _T_5117_33; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_449 = _T_4843 ? _T_4292_34 : _T_5117_34; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_450 = _T_4843 ? _T_4292_35 : _T_5117_35; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_451 = _T_4843 ? _T_4292_36 : _T_5117_36; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_452 = _T_4843 ? _T_4292_37 : _T_5117_37; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_453 = _T_4843 ? _T_4292_38 : _T_5117_38; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_454 = _T_4843 ? _T_4292_39 : _T_5117_39; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_455 = _T_4843 ? _T_4292_40 : _T_5117_40; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_456 = _T_4843 ? _T_4292_41 : _T_5117_41; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_457 = _T_4843 ? _T_4292_42 : _T_5117_42; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_458 = _T_4843 ? _T_4292_43 : _T_5117_43; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_459 = _T_4843 ? _T_4292_44 : _T_5117_44; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_460 = _T_4843 ? _T_4292_45 : _T_5117_45; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_461 = _T_4843 ? _T_4292_46 : _T_5117_46; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_462 = _T_4843 ? _T_4292_47 : _T_5117_47; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_463 = _T_4843 ? _T_4292_48 : _T_5117_48; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_464 = _T_4843 ? _T_4292_49 : _T_5117_49; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_465 = _T_4843 ? _T_4292_50 : _T_5117_50; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_466 = _T_4843 ? _T_4292_51 : _T_5117_51; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_467 = _T_4843 ? _T_4292_52 : _T_5117_52; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_468 = _T_4843 ? _T_4292_53 : _T_5117_53; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_469 = _T_4843 ? _T_4292_54 : _T_5117_54; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_470 = _T_4843 ? _T_4292_55 : _T_5117_55; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_471 = _T_4843 ? _T_4292_56 : _T_5117_56; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_472 = _T_4843 ? _T_4292_57 : _T_5117_57; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_473 = _T_4843 ? _T_4292_58 : _T_5117_58; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_474 = _T_4843 ? _T_4292_59 : _T_5117_59; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_475 = _T_4843 ? _T_4292_60 : _T_5117_60; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_476 = _T_4843 ? _T_4292_61 : _T_5117_61; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_477 = _T_4843 ? _T_4292_62 : _T_5117_62; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_478 = _T_4843 ? _T_4292_63 : _T_5117_63; // @[Reg.scala 20:19:@3012.4]
  assign _GEN_479 = _T_4843 ? _T_4292_0 : _T_5581_0; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_480 = _T_4843 ? _T_4292_1 : _T_5581_1; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_481 = _T_4843 ? _T_4292_2 : _T_5581_2; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_482 = _T_4843 ? _T_4292_3 : _T_5581_3; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_483 = _T_4843 ? _T_4292_4 : _T_5581_4; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_484 = _T_4843 ? _T_4292_5 : _T_5581_5; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_485 = _T_4843 ? _T_4292_6 : _T_5581_6; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_486 = _T_4843 ? _T_4292_7 : _T_5581_7; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_487 = _T_4843 ? _T_4292_8 : _T_5581_8; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_488 = _T_4843 ? _T_4292_9 : _T_5581_9; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_489 = _T_4843 ? _T_4292_10 : _T_5581_10; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_490 = _T_4843 ? _T_4292_11 : _T_5581_11; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_491 = _T_4843 ? _T_4292_12 : _T_5581_12; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_492 = _T_4843 ? _T_4292_13 : _T_5581_13; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_493 = _T_4843 ? _T_4292_14 : _T_5581_14; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_494 = _T_4843 ? _T_4292_15 : _T_5581_15; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_495 = _T_4843 ? _T_4292_16 : _T_5581_16; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_496 = _T_4843 ? _T_4292_17 : _T_5581_17; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_497 = _T_4843 ? _T_4292_18 : _T_5581_18; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_498 = _T_4843 ? _T_4292_19 : _T_5581_19; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_499 = _T_4843 ? _T_4292_20 : _T_5581_20; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_500 = _T_4843 ? _T_4292_21 : _T_5581_21; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_501 = _T_4843 ? _T_4292_22 : _T_5581_22; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_502 = _T_4843 ? _T_4292_23 : _T_5581_23; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_503 = _T_4843 ? _T_4292_24 : _T_5581_24; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_504 = _T_4843 ? _T_4292_25 : _T_5581_25; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_505 = _T_4843 ? _T_4292_26 : _T_5581_26; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_506 = _T_4843 ? _T_4292_27 : _T_5581_27; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_507 = _T_4843 ? _T_4292_28 : _T_5581_28; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_508 = _T_4843 ? _T_4292_29 : _T_5581_29; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_509 = _T_4843 ? _T_4292_30 : _T_5581_30; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_510 = _T_4843 ? _T_4292_31 : _T_5581_31; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_511 = _T_4843 ? _T_4292_32 : _T_5581_32; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_512 = _T_4843 ? _T_4292_33 : _T_5581_33; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_513 = _T_4843 ? _T_4292_34 : _T_5581_34; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_514 = _T_4843 ? _T_4292_35 : _T_5581_35; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_515 = _T_4843 ? _T_4292_36 : _T_5581_36; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_516 = _T_4843 ? _T_4292_37 : _T_5581_37; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_517 = _T_4843 ? _T_4292_38 : _T_5581_38; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_518 = _T_4843 ? _T_4292_39 : _T_5581_39; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_519 = _T_4843 ? _T_4292_40 : _T_5581_40; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_520 = _T_4843 ? _T_4292_41 : _T_5581_41; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_521 = _T_4843 ? _T_4292_42 : _T_5581_42; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_522 = _T_4843 ? _T_4292_43 : _T_5581_43; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_523 = _T_4843 ? _T_4292_44 : _T_5581_44; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_524 = _T_4843 ? _T_4292_45 : _T_5581_45; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_525 = _T_4843 ? _T_4292_46 : _T_5581_46; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_526 = _T_4843 ? _T_4292_47 : _T_5581_47; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_527 = _T_4843 ? _T_4292_48 : _T_5581_48; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_528 = _T_4843 ? _T_4292_49 : _T_5581_49; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_529 = _T_4843 ? _T_4292_50 : _T_5581_50; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_530 = _T_4843 ? _T_4292_51 : _T_5581_51; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_531 = _T_4843 ? _T_4292_52 : _T_5581_52; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_532 = _T_4843 ? _T_4292_53 : _T_5581_53; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_533 = _T_4843 ? _T_4292_54 : _T_5581_54; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_534 = _T_4843 ? _T_4292_55 : _T_5581_55; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_535 = _T_4843 ? _T_4292_56 : _T_5581_56; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_536 = _T_4843 ? _T_4292_57 : _T_5581_57; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_537 = _T_4843 ? _T_4292_58 : _T_5581_58; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_538 = _T_4843 ? _T_4292_59 : _T_5581_59; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_539 = _T_4843 ? _T_4292_60 : _T_5581_60; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_540 = _T_4843 ? _T_4292_61 : _T_5581_61; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_541 = _T_4843 ? _T_4292_62 : _T_5581_62; // @[Reg.scala 20:19:@3209.4]
  assign _GEN_542 = _T_4843 ? _T_4292_63 : _T_5581_63; // @[Reg.scala 20:19:@3209.4]
  assign io_sc2cdma_dat_updt_valid = _T_1169; // @[NV_NVDLA_CSC_dl_for_check.scala 310:27:@326.4]
  assign io_sc2cdma_dat_updt_bits_entries = _T_1175; // @[NV_NVDLA_CSC_dl_for_check.scala 312:34:@336.4]
  assign io_sc2cdma_dat_updt_bits_slices = _T_1172; // @[NV_NVDLA_CSC_dl_for_check.scala 311:33:@331.4]
  assign io_sc2buf_dat_rd_addr_valid = _T_1781; // @[NV_NVDLA_CSC_dl_for_check.scala 727:29:@933.4]
  assign io_sc2buf_dat_rd_addr_bits = _T_1788[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 728:28:@934.4]
  assign io_sc2mac_dat_a_valid = _T_4838; // @[NV_NVDLA_CSC_dl_for_check.scala 1176:23:@2929.4]
  assign io_sc2mac_dat_a_bits_mask_0 = _T_5117_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3078.4]
  assign io_sc2mac_dat_a_bits_mask_1 = _T_5117_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3079.4]
  assign io_sc2mac_dat_a_bits_mask_2 = _T_5117_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3080.4]
  assign io_sc2mac_dat_a_bits_mask_3 = _T_5117_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3081.4]
  assign io_sc2mac_dat_a_bits_mask_4 = _T_5117_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3082.4]
  assign io_sc2mac_dat_a_bits_mask_5 = _T_5117_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3083.4]
  assign io_sc2mac_dat_a_bits_mask_6 = _T_5117_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3084.4]
  assign io_sc2mac_dat_a_bits_mask_7 = _T_5117_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3085.4]
  assign io_sc2mac_dat_a_bits_mask_8 = _T_5117_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3086.4]
  assign io_sc2mac_dat_a_bits_mask_9 = _T_5117_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3087.4]
  assign io_sc2mac_dat_a_bits_mask_10 = _T_5117_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3088.4]
  assign io_sc2mac_dat_a_bits_mask_11 = _T_5117_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3089.4]
  assign io_sc2mac_dat_a_bits_mask_12 = _T_5117_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3090.4]
  assign io_sc2mac_dat_a_bits_mask_13 = _T_5117_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3091.4]
  assign io_sc2mac_dat_a_bits_mask_14 = _T_5117_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3092.4]
  assign io_sc2mac_dat_a_bits_mask_15 = _T_5117_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3093.4]
  assign io_sc2mac_dat_a_bits_mask_16 = _T_5117_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3094.4]
  assign io_sc2mac_dat_a_bits_mask_17 = _T_5117_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3095.4]
  assign io_sc2mac_dat_a_bits_mask_18 = _T_5117_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3096.4]
  assign io_sc2mac_dat_a_bits_mask_19 = _T_5117_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3097.4]
  assign io_sc2mac_dat_a_bits_mask_20 = _T_5117_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3098.4]
  assign io_sc2mac_dat_a_bits_mask_21 = _T_5117_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3099.4]
  assign io_sc2mac_dat_a_bits_mask_22 = _T_5117_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3100.4]
  assign io_sc2mac_dat_a_bits_mask_23 = _T_5117_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3101.4]
  assign io_sc2mac_dat_a_bits_mask_24 = _T_5117_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3102.4]
  assign io_sc2mac_dat_a_bits_mask_25 = _T_5117_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3103.4]
  assign io_sc2mac_dat_a_bits_mask_26 = _T_5117_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3104.4]
  assign io_sc2mac_dat_a_bits_mask_27 = _T_5117_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3105.4]
  assign io_sc2mac_dat_a_bits_mask_28 = _T_5117_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3106.4]
  assign io_sc2mac_dat_a_bits_mask_29 = _T_5117_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3107.4]
  assign io_sc2mac_dat_a_bits_mask_30 = _T_5117_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3108.4]
  assign io_sc2mac_dat_a_bits_mask_31 = _T_5117_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3109.4]
  assign io_sc2mac_dat_a_bits_mask_32 = _T_5117_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3110.4]
  assign io_sc2mac_dat_a_bits_mask_33 = _T_5117_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3111.4]
  assign io_sc2mac_dat_a_bits_mask_34 = _T_5117_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3112.4]
  assign io_sc2mac_dat_a_bits_mask_35 = _T_5117_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3113.4]
  assign io_sc2mac_dat_a_bits_mask_36 = _T_5117_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3114.4]
  assign io_sc2mac_dat_a_bits_mask_37 = _T_5117_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3115.4]
  assign io_sc2mac_dat_a_bits_mask_38 = _T_5117_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3116.4]
  assign io_sc2mac_dat_a_bits_mask_39 = _T_5117_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3117.4]
  assign io_sc2mac_dat_a_bits_mask_40 = _T_5117_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3118.4]
  assign io_sc2mac_dat_a_bits_mask_41 = _T_5117_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3119.4]
  assign io_sc2mac_dat_a_bits_mask_42 = _T_5117_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3120.4]
  assign io_sc2mac_dat_a_bits_mask_43 = _T_5117_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3121.4]
  assign io_sc2mac_dat_a_bits_mask_44 = _T_5117_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3122.4]
  assign io_sc2mac_dat_a_bits_mask_45 = _T_5117_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3123.4]
  assign io_sc2mac_dat_a_bits_mask_46 = _T_5117_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3124.4]
  assign io_sc2mac_dat_a_bits_mask_47 = _T_5117_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3125.4]
  assign io_sc2mac_dat_a_bits_mask_48 = _T_5117_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3126.4]
  assign io_sc2mac_dat_a_bits_mask_49 = _T_5117_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3127.4]
  assign io_sc2mac_dat_a_bits_mask_50 = _T_5117_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3128.4]
  assign io_sc2mac_dat_a_bits_mask_51 = _T_5117_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3129.4]
  assign io_sc2mac_dat_a_bits_mask_52 = _T_5117_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3130.4]
  assign io_sc2mac_dat_a_bits_mask_53 = _T_5117_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3131.4]
  assign io_sc2mac_dat_a_bits_mask_54 = _T_5117_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3132.4]
  assign io_sc2mac_dat_a_bits_mask_55 = _T_5117_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3133.4]
  assign io_sc2mac_dat_a_bits_mask_56 = _T_5117_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3134.4]
  assign io_sc2mac_dat_a_bits_mask_57 = _T_5117_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3135.4]
  assign io_sc2mac_dat_a_bits_mask_58 = _T_5117_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3136.4]
  assign io_sc2mac_dat_a_bits_mask_59 = _T_5117_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3137.4]
  assign io_sc2mac_dat_a_bits_mask_60 = _T_5117_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3138.4]
  assign io_sc2mac_dat_a_bits_mask_61 = _T_5117_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3139.4]
  assign io_sc2mac_dat_a_bits_mask_62 = _T_5117_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3140.4]
  assign io_sc2mac_dat_a_bits_mask_63 = _T_5117_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1180:27:@3141.4]
  assign io_sc2mac_dat_a_bits_data_0 = _T_5779; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3343.4]
  assign io_sc2mac_dat_a_bits_data_1 = _T_5783; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3353.4]
  assign io_sc2mac_dat_a_bits_data_2 = _T_5787; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3363.4]
  assign io_sc2mac_dat_a_bits_data_3 = _T_5791; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3373.4]
  assign io_sc2mac_dat_a_bits_data_4 = _T_5795; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3383.4]
  assign io_sc2mac_dat_a_bits_data_5 = _T_5799; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3393.4]
  assign io_sc2mac_dat_a_bits_data_6 = _T_5803; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3403.4]
  assign io_sc2mac_dat_a_bits_data_7 = _T_5807; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3413.4]
  assign io_sc2mac_dat_a_bits_data_8 = _T_5811; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3423.4]
  assign io_sc2mac_dat_a_bits_data_9 = _T_5815; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3433.4]
  assign io_sc2mac_dat_a_bits_data_10 = _T_5819; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3443.4]
  assign io_sc2mac_dat_a_bits_data_11 = _T_5823; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3453.4]
  assign io_sc2mac_dat_a_bits_data_12 = _T_5827; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3463.4]
  assign io_sc2mac_dat_a_bits_data_13 = _T_5831; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3473.4]
  assign io_sc2mac_dat_a_bits_data_14 = _T_5835; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3483.4]
  assign io_sc2mac_dat_a_bits_data_15 = _T_5839; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3493.4]
  assign io_sc2mac_dat_a_bits_data_16 = _T_5843; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3503.4]
  assign io_sc2mac_dat_a_bits_data_17 = _T_5847; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3513.4]
  assign io_sc2mac_dat_a_bits_data_18 = _T_5851; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3523.4]
  assign io_sc2mac_dat_a_bits_data_19 = _T_5855; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3533.4]
  assign io_sc2mac_dat_a_bits_data_20 = _T_5859; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3543.4]
  assign io_sc2mac_dat_a_bits_data_21 = _T_5863; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3553.4]
  assign io_sc2mac_dat_a_bits_data_22 = _T_5867; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3563.4]
  assign io_sc2mac_dat_a_bits_data_23 = _T_5871; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3573.4]
  assign io_sc2mac_dat_a_bits_data_24 = _T_5875; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3583.4]
  assign io_sc2mac_dat_a_bits_data_25 = _T_5879; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3593.4]
  assign io_sc2mac_dat_a_bits_data_26 = _T_5883; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3603.4]
  assign io_sc2mac_dat_a_bits_data_27 = _T_5887; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3613.4]
  assign io_sc2mac_dat_a_bits_data_28 = _T_5891; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3623.4]
  assign io_sc2mac_dat_a_bits_data_29 = _T_5895; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3633.4]
  assign io_sc2mac_dat_a_bits_data_30 = _T_5899; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3643.4]
  assign io_sc2mac_dat_a_bits_data_31 = _T_5903; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3653.4]
  assign io_sc2mac_dat_a_bits_data_32 = _T_5907; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3663.4]
  assign io_sc2mac_dat_a_bits_data_33 = _T_5911; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3673.4]
  assign io_sc2mac_dat_a_bits_data_34 = _T_5915; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3683.4]
  assign io_sc2mac_dat_a_bits_data_35 = _T_5919; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3693.4]
  assign io_sc2mac_dat_a_bits_data_36 = _T_5923; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3703.4]
  assign io_sc2mac_dat_a_bits_data_37 = _T_5927; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3713.4]
  assign io_sc2mac_dat_a_bits_data_38 = _T_5931; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3723.4]
  assign io_sc2mac_dat_a_bits_data_39 = _T_5935; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3733.4]
  assign io_sc2mac_dat_a_bits_data_40 = _T_5939; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3743.4]
  assign io_sc2mac_dat_a_bits_data_41 = _T_5943; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3753.4]
  assign io_sc2mac_dat_a_bits_data_42 = _T_5947; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3763.4]
  assign io_sc2mac_dat_a_bits_data_43 = _T_5951; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3773.4]
  assign io_sc2mac_dat_a_bits_data_44 = _T_5955; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3783.4]
  assign io_sc2mac_dat_a_bits_data_45 = _T_5959; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3793.4]
  assign io_sc2mac_dat_a_bits_data_46 = _T_5963; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3803.4]
  assign io_sc2mac_dat_a_bits_data_47 = _T_5967; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3813.4]
  assign io_sc2mac_dat_a_bits_data_48 = _T_5971; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3823.4]
  assign io_sc2mac_dat_a_bits_data_49 = _T_5975; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3833.4]
  assign io_sc2mac_dat_a_bits_data_50 = _T_5979; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3843.4]
  assign io_sc2mac_dat_a_bits_data_51 = _T_5983; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3853.4]
  assign io_sc2mac_dat_a_bits_data_52 = _T_5987; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3863.4]
  assign io_sc2mac_dat_a_bits_data_53 = _T_5991; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3873.4]
  assign io_sc2mac_dat_a_bits_data_54 = _T_5995; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3883.4]
  assign io_sc2mac_dat_a_bits_data_55 = _T_5999; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3893.4]
  assign io_sc2mac_dat_a_bits_data_56 = _T_6003; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3903.4]
  assign io_sc2mac_dat_a_bits_data_57 = _T_6007; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3913.4]
  assign io_sc2mac_dat_a_bits_data_58 = _T_6011; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3923.4]
  assign io_sc2mac_dat_a_bits_data_59 = _T_6015; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3933.4]
  assign io_sc2mac_dat_a_bits_data_60 = _T_6019; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3943.4]
  assign io_sc2mac_dat_a_bits_data_61 = _T_6023; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3953.4]
  assign io_sc2mac_dat_a_bits_data_62 = _T_6027; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3963.4]
  assign io_sc2mac_dat_a_bits_data_63 = _T_6031; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:34:@3973.4]
  assign io_sc2mac_dat_a_bits_pd = _T_4845; // @[NV_NVDLA_CSC_dl_for_check.scala 1178:25:@2938.4]
  assign io_sc2mac_dat_b_valid = _T_4841; // @[NV_NVDLA_CSC_dl_for_check.scala 1177:23:@2932.4]
  assign io_sc2mac_dat_b_bits_mask_0 = _T_5581_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3275.4]
  assign io_sc2mac_dat_b_bits_mask_1 = _T_5581_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3276.4]
  assign io_sc2mac_dat_b_bits_mask_2 = _T_5581_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3277.4]
  assign io_sc2mac_dat_b_bits_mask_3 = _T_5581_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3278.4]
  assign io_sc2mac_dat_b_bits_mask_4 = _T_5581_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3279.4]
  assign io_sc2mac_dat_b_bits_mask_5 = _T_5581_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3280.4]
  assign io_sc2mac_dat_b_bits_mask_6 = _T_5581_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3281.4]
  assign io_sc2mac_dat_b_bits_mask_7 = _T_5581_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3282.4]
  assign io_sc2mac_dat_b_bits_mask_8 = _T_5581_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3283.4]
  assign io_sc2mac_dat_b_bits_mask_9 = _T_5581_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3284.4]
  assign io_sc2mac_dat_b_bits_mask_10 = _T_5581_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3285.4]
  assign io_sc2mac_dat_b_bits_mask_11 = _T_5581_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3286.4]
  assign io_sc2mac_dat_b_bits_mask_12 = _T_5581_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3287.4]
  assign io_sc2mac_dat_b_bits_mask_13 = _T_5581_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3288.4]
  assign io_sc2mac_dat_b_bits_mask_14 = _T_5581_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3289.4]
  assign io_sc2mac_dat_b_bits_mask_15 = _T_5581_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3290.4]
  assign io_sc2mac_dat_b_bits_mask_16 = _T_5581_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3291.4]
  assign io_sc2mac_dat_b_bits_mask_17 = _T_5581_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3292.4]
  assign io_sc2mac_dat_b_bits_mask_18 = _T_5581_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3293.4]
  assign io_sc2mac_dat_b_bits_mask_19 = _T_5581_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3294.4]
  assign io_sc2mac_dat_b_bits_mask_20 = _T_5581_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3295.4]
  assign io_sc2mac_dat_b_bits_mask_21 = _T_5581_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3296.4]
  assign io_sc2mac_dat_b_bits_mask_22 = _T_5581_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3297.4]
  assign io_sc2mac_dat_b_bits_mask_23 = _T_5581_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3298.4]
  assign io_sc2mac_dat_b_bits_mask_24 = _T_5581_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3299.4]
  assign io_sc2mac_dat_b_bits_mask_25 = _T_5581_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3300.4]
  assign io_sc2mac_dat_b_bits_mask_26 = _T_5581_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3301.4]
  assign io_sc2mac_dat_b_bits_mask_27 = _T_5581_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3302.4]
  assign io_sc2mac_dat_b_bits_mask_28 = _T_5581_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3303.4]
  assign io_sc2mac_dat_b_bits_mask_29 = _T_5581_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3304.4]
  assign io_sc2mac_dat_b_bits_mask_30 = _T_5581_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3305.4]
  assign io_sc2mac_dat_b_bits_mask_31 = _T_5581_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3306.4]
  assign io_sc2mac_dat_b_bits_mask_32 = _T_5581_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3307.4]
  assign io_sc2mac_dat_b_bits_mask_33 = _T_5581_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3308.4]
  assign io_sc2mac_dat_b_bits_mask_34 = _T_5581_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3309.4]
  assign io_sc2mac_dat_b_bits_mask_35 = _T_5581_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3310.4]
  assign io_sc2mac_dat_b_bits_mask_36 = _T_5581_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3311.4]
  assign io_sc2mac_dat_b_bits_mask_37 = _T_5581_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3312.4]
  assign io_sc2mac_dat_b_bits_mask_38 = _T_5581_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3313.4]
  assign io_sc2mac_dat_b_bits_mask_39 = _T_5581_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3314.4]
  assign io_sc2mac_dat_b_bits_mask_40 = _T_5581_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3315.4]
  assign io_sc2mac_dat_b_bits_mask_41 = _T_5581_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3316.4]
  assign io_sc2mac_dat_b_bits_mask_42 = _T_5581_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3317.4]
  assign io_sc2mac_dat_b_bits_mask_43 = _T_5581_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3318.4]
  assign io_sc2mac_dat_b_bits_mask_44 = _T_5581_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3319.4]
  assign io_sc2mac_dat_b_bits_mask_45 = _T_5581_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3320.4]
  assign io_sc2mac_dat_b_bits_mask_46 = _T_5581_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3321.4]
  assign io_sc2mac_dat_b_bits_mask_47 = _T_5581_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3322.4]
  assign io_sc2mac_dat_b_bits_mask_48 = _T_5581_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3323.4]
  assign io_sc2mac_dat_b_bits_mask_49 = _T_5581_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3324.4]
  assign io_sc2mac_dat_b_bits_mask_50 = _T_5581_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3325.4]
  assign io_sc2mac_dat_b_bits_mask_51 = _T_5581_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3326.4]
  assign io_sc2mac_dat_b_bits_mask_52 = _T_5581_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3327.4]
  assign io_sc2mac_dat_b_bits_mask_53 = _T_5581_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3328.4]
  assign io_sc2mac_dat_b_bits_mask_54 = _T_5581_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3329.4]
  assign io_sc2mac_dat_b_bits_mask_55 = _T_5581_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3330.4]
  assign io_sc2mac_dat_b_bits_mask_56 = _T_5581_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3331.4]
  assign io_sc2mac_dat_b_bits_mask_57 = _T_5581_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3332.4]
  assign io_sc2mac_dat_b_bits_mask_58 = _T_5581_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3333.4]
  assign io_sc2mac_dat_b_bits_mask_59 = _T_5581_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3334.4]
  assign io_sc2mac_dat_b_bits_mask_60 = _T_5581_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3335.4]
  assign io_sc2mac_dat_b_bits_mask_61 = _T_5581_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3336.4]
  assign io_sc2mac_dat_b_bits_mask_62 = _T_5581_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3337.4]
  assign io_sc2mac_dat_b_bits_mask_63 = _T_5581_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1181:27:@3338.4]
  assign io_sc2mac_dat_b_bits_data_0 = _T_5781; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3348.4]
  assign io_sc2mac_dat_b_bits_data_1 = _T_5785; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3358.4]
  assign io_sc2mac_dat_b_bits_data_2 = _T_5789; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3368.4]
  assign io_sc2mac_dat_b_bits_data_3 = _T_5793; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3378.4]
  assign io_sc2mac_dat_b_bits_data_4 = _T_5797; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3388.4]
  assign io_sc2mac_dat_b_bits_data_5 = _T_5801; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3398.4]
  assign io_sc2mac_dat_b_bits_data_6 = _T_5805; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3408.4]
  assign io_sc2mac_dat_b_bits_data_7 = _T_5809; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3418.4]
  assign io_sc2mac_dat_b_bits_data_8 = _T_5813; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3428.4]
  assign io_sc2mac_dat_b_bits_data_9 = _T_5817; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3438.4]
  assign io_sc2mac_dat_b_bits_data_10 = _T_5821; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3448.4]
  assign io_sc2mac_dat_b_bits_data_11 = _T_5825; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3458.4]
  assign io_sc2mac_dat_b_bits_data_12 = _T_5829; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3468.4]
  assign io_sc2mac_dat_b_bits_data_13 = _T_5833; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3478.4]
  assign io_sc2mac_dat_b_bits_data_14 = _T_5837; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3488.4]
  assign io_sc2mac_dat_b_bits_data_15 = _T_5841; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3498.4]
  assign io_sc2mac_dat_b_bits_data_16 = _T_5845; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3508.4]
  assign io_sc2mac_dat_b_bits_data_17 = _T_5849; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3518.4]
  assign io_sc2mac_dat_b_bits_data_18 = _T_5853; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3528.4]
  assign io_sc2mac_dat_b_bits_data_19 = _T_5857; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3538.4]
  assign io_sc2mac_dat_b_bits_data_20 = _T_5861; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3548.4]
  assign io_sc2mac_dat_b_bits_data_21 = _T_5865; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3558.4]
  assign io_sc2mac_dat_b_bits_data_22 = _T_5869; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3568.4]
  assign io_sc2mac_dat_b_bits_data_23 = _T_5873; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3578.4]
  assign io_sc2mac_dat_b_bits_data_24 = _T_5877; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3588.4]
  assign io_sc2mac_dat_b_bits_data_25 = _T_5881; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3598.4]
  assign io_sc2mac_dat_b_bits_data_26 = _T_5885; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3608.4]
  assign io_sc2mac_dat_b_bits_data_27 = _T_5889; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3618.4]
  assign io_sc2mac_dat_b_bits_data_28 = _T_5893; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3628.4]
  assign io_sc2mac_dat_b_bits_data_29 = _T_5897; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3638.4]
  assign io_sc2mac_dat_b_bits_data_30 = _T_5901; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3648.4]
  assign io_sc2mac_dat_b_bits_data_31 = _T_5905; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3658.4]
  assign io_sc2mac_dat_b_bits_data_32 = _T_5909; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3668.4]
  assign io_sc2mac_dat_b_bits_data_33 = _T_5913; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3678.4]
  assign io_sc2mac_dat_b_bits_data_34 = _T_5917; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3688.4]
  assign io_sc2mac_dat_b_bits_data_35 = _T_5921; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3698.4]
  assign io_sc2mac_dat_b_bits_data_36 = _T_5925; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3708.4]
  assign io_sc2mac_dat_b_bits_data_37 = _T_5929; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3718.4]
  assign io_sc2mac_dat_b_bits_data_38 = _T_5933; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3728.4]
  assign io_sc2mac_dat_b_bits_data_39 = _T_5937; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3738.4]
  assign io_sc2mac_dat_b_bits_data_40 = _T_5941; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3748.4]
  assign io_sc2mac_dat_b_bits_data_41 = _T_5945; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3758.4]
  assign io_sc2mac_dat_b_bits_data_42 = _T_5949; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3768.4]
  assign io_sc2mac_dat_b_bits_data_43 = _T_5953; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3778.4]
  assign io_sc2mac_dat_b_bits_data_44 = _T_5957; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3788.4]
  assign io_sc2mac_dat_b_bits_data_45 = _T_5961; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3798.4]
  assign io_sc2mac_dat_b_bits_data_46 = _T_5965; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3808.4]
  assign io_sc2mac_dat_b_bits_data_47 = _T_5969; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3818.4]
  assign io_sc2mac_dat_b_bits_data_48 = _T_5973; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3828.4]
  assign io_sc2mac_dat_b_bits_data_49 = _T_5977; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3838.4]
  assign io_sc2mac_dat_b_bits_data_50 = _T_5981; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3848.4]
  assign io_sc2mac_dat_b_bits_data_51 = _T_5985; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3858.4]
  assign io_sc2mac_dat_b_bits_data_52 = _T_5989; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3868.4]
  assign io_sc2mac_dat_b_bits_data_53 = _T_5993; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3878.4]
  assign io_sc2mac_dat_b_bits_data_54 = _T_5997; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3888.4]
  assign io_sc2mac_dat_b_bits_data_55 = _T_6001; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3898.4]
  assign io_sc2mac_dat_b_bits_data_56 = _T_6005; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3908.4]
  assign io_sc2mac_dat_b_bits_data_57 = _T_6009; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3918.4]
  assign io_sc2mac_dat_b_bits_data_58 = _T_6013; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3928.4]
  assign io_sc2mac_dat_b_bits_data_59 = _T_6017; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3938.4]
  assign io_sc2mac_dat_b_bits_data_60 = _T_6021; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3948.4]
  assign io_sc2mac_dat_b_bits_data_61 = _T_6025; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3958.4]
  assign io_sc2mac_dat_b_bits_data_62 = _T_6029; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3968.4]
  assign io_sc2mac_dat_b_bits_data_63 = _T_6033; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:34:@3978.4]
  assign io_sc2mac_dat_b_bits_pd = _T_4849; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:25:@2944.4]
  assign io_slcg_wg_en = 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 251:15:@243.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_718 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_725 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_732 = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_739 = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_746 = _RAND_4[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_753 = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_760 = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_774 = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_781 = _RAND_8[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_788 = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_795 = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  _T_834 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_841 = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_848 = _RAND_13[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_855 = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_862 = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_869 = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_872 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_875 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_881 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_884 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_887 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_890 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_896 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_899 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_905 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_908 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_911 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_918 = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_925 = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_935 = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_942 = _RAND_31[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_949 = _RAND_32[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_956 = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_963 = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_970 = _RAND_35[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_977 = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_984 = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_991 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_998 = _RAND_39[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_1005 = _RAND_40[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_1012 = _RAND_41[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_1019 = _RAND_42[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_1026 = _RAND_43[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_1079 = _RAND_44[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_2220 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_2214 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_2211 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_2234 = _RAND_48[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_2228 = _RAND_49[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_2225 = _RAND_50[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1169 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1172 = _RAND_52[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_1175 = _RAND_53[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_1180 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_1183 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_1186 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_1189 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_1192 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_1214 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_1217 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_1220 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_1223 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_1228 = _RAND_63[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_1231 = _RAND_64[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_1234 = _RAND_65[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_1237 = _RAND_66[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_1282 = _RAND_67[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_1293 = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_1309 = _RAND_69[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_1338 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_1332 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_1335 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_1364 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_1369 = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_1372 = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1393 = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1407 = _RAND_77[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_1410 = _RAND_78[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_1413 = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_1416 = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_1419 = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_1422 = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_1427 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_1430 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_1542 = _RAND_85[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_1545 = _RAND_86[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_1619 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_1622 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_1625 = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_1628 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_1631 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_1634 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_1637 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_1640 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_1643 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_1646 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_1651 = _RAND_97[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_1654 = _RAND_98[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_1657 = _RAND_99[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_1660 = _RAND_100[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_1663 = _RAND_101[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_1666 = _RAND_102[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_1669 = _RAND_103[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_1762_0 = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_1762_1 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_1762_2 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_1762_3 = _RAND_107[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_1781 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_1788 = _RAND_109[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_1791 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_1797 = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_1800 = _RAND_112[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_1803 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_1806 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_1809 = _RAND_115[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_1812 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_1815 = _RAND_117[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_1818 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_1821 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1824 = _RAND_120[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1946 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1949 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1952 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1955 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_1958 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1961 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1966 = _RAND_127[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1969 = _RAND_128[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1972 = _RAND_129[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1975 = _RAND_130[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1978 = _RAND_131[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1981 = _RAND_132[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_2054 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_2066 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {16{`RANDOM}};
  _T_2077 = _RAND_135[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {16{`RANDOM}};
  _T_2085 = _RAND_136[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_2185 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_2188 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_2191 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_2194 = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_2197 = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_2200 = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_2203 = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_2206 = _RAND_144[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_2217 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_2231 = _RAND_146[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {8{`RANDOM}};
  _T_2614 = _RAND_147[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {4{`RANDOM}};
  _T_2616 = _RAND_148[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {4{`RANDOM}};
  _T_2618 = _RAND_149[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {4{`RANDOM}};
  _T_2620 = _RAND_150[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {4{`RANDOM}};
  _T_2622 = _RAND_151[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {4{`RANDOM}};
  _T_2624 = _RAND_152[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_3422 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_3692_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_3692_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_3692_2 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_3692_3 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_3692_4 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_3692_5 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_3692_6 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_3692_7 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_3692_8 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_3692_9 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_3692_10 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_3692_11 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_3692_12 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_3692_13 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_3692_14 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_3692_15 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_3692_16 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_3692_17 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_3692_18 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_3692_19 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_3692_20 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_3692_21 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_3692_22 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_3692_23 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_3692_24 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_3692_25 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_3692_26 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_3692_27 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_3692_28 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_3692_29 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_3692_30 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_3692_31 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_3692_32 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_3692_33 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_3692_34 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_3692_35 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_3692_36 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_3692_37 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_3692_38 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_3692_39 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_3692_40 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_3692_41 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_3692_42 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_3692_43 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_3692_44 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_3692_45 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_3692_46 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_3692_47 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_3692_48 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_3692_49 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_3692_50 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_3692_51 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_3692_52 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_3692_53 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_3692_54 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_3692_55 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_3692_56 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_3692_57 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_3692_58 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_3692_59 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_3692_60 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_3692_61 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_3692_62 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_3692_63 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_3892_0 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_3892_1 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_3892_2 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_3892_3 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_3892_4 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_3892_5 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_3892_6 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_3892_7 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_3892_8 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_3892_9 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_3892_10 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_3892_11 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_3892_12 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_3892_13 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_3892_14 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_3892_15 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_3892_16 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_3892_17 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_3892_18 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_3892_19 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_3892_20 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_3892_21 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_3892_22 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_3892_23 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_3892_24 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_3892_25 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_3892_26 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_3892_27 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_3892_28 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_3892_29 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_3892_30 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_3892_31 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_3892_32 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_3892_33 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_3892_34 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_3892_35 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_3892_36 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_3892_37 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_3892_38 = _RAND_256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_3892_39 = _RAND_257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_3892_40 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_3892_41 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_3892_42 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_3892_43 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_3892_44 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_3892_45 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_3892_46 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_3892_47 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_3892_48 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_3892_49 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_3892_50 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_3892_51 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_3892_52 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_3892_53 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_3892_54 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_3892_55 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_3892_56 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_3892_57 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_3892_58 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_3892_59 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_3892_60 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_3892_61 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_3892_62 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_3892_63 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_4025 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_4292_0 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_4292_1 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_4292_2 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_4292_3 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_4292_4 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_4292_5 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_4292_6 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_4292_7 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_4292_8 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_4292_9 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_4292_10 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_4292_11 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_4292_12 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_4292_13 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_4292_14 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_4292_15 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_4292_16 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_4292_17 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_4292_18 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_4292_19 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_4292_20 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_4292_21 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_4292_22 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_4292_23 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_4292_24 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_4292_25 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_4292_26 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_4292_27 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_4292_28 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_4292_29 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_4292_30 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_4292_31 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_4292_32 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_4292_33 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_4292_34 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_4292_35 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_4292_36 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_4292_37 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_4292_38 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_4292_39 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_4292_40 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_4292_41 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_4292_42 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_4292_43 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_4292_44 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_4292_45 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_4292_46 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_4292_47 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_4292_48 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_4292_49 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_4292_50 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_4292_51 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_4292_52 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_4292_53 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_4292_54 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_4292_55 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_4292_56 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_4292_57 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_4292_58 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_4292_59 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_4292_60 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_4292_61 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_4292_62 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_4292_63 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_4491 = _RAND_347[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_4495_0 = _RAND_348[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_4495_1 = _RAND_349[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_4495_2 = _RAND_350[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_4495_3 = _RAND_351[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_4495_4 = _RAND_352[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_4495_5 = _RAND_353[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_4495_6 = _RAND_354[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_4495_7 = _RAND_355[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_4495_8 = _RAND_356[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_4495_9 = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_4495_10 = _RAND_358[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_4495_11 = _RAND_359[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_4495_12 = _RAND_360[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_4495_13 = _RAND_361[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_4495_14 = _RAND_362[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_4495_15 = _RAND_363[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_4495_16 = _RAND_364[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_4495_17 = _RAND_365[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_4495_18 = _RAND_366[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_4495_19 = _RAND_367[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_4495_20 = _RAND_368[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_4495_21 = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_4495_22 = _RAND_370[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_4495_23 = _RAND_371[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_4495_24 = _RAND_372[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_4495_25 = _RAND_373[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_4495_26 = _RAND_374[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_4495_27 = _RAND_375[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_4495_28 = _RAND_376[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_4495_29 = _RAND_377[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_4495_30 = _RAND_378[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_4495_31 = _RAND_379[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_4495_32 = _RAND_380[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_4495_33 = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_4495_34 = _RAND_382[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_4495_35 = _RAND_383[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_4495_36 = _RAND_384[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_4495_37 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_4495_38 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_4495_39 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_4495_40 = _RAND_388[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_4495_41 = _RAND_389[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_4495_42 = _RAND_390[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_4495_43 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_4495_44 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_4495_45 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_4495_46 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_4495_47 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_4495_48 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_4495_49 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_4495_50 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_4495_51 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_4495_52 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_4495_53 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_4495_54 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_4495_55 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_4495_56 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_4495_57 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_4495_58 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_4495_59 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_4495_60 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_4495_61 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_4495_62 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_4495_63 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_4832 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4838 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4841 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4845 = _RAND_415[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4849 = _RAND_416[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_5117_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_5117_1 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_5117_2 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_5117_3 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_5117_4 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_5117_5 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_5117_6 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_5117_7 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_5117_8 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_5117_9 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_5117_10 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_5117_11 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_5117_12 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_5117_13 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_5117_14 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_5117_15 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_5117_16 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_5117_17 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_5117_18 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_5117_19 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_5117_20 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_5117_21 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_5117_22 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_5117_23 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_5117_24 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_5117_25 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_5117_26 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_5117_27 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_5117_28 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_5117_29 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_5117_30 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_5117_31 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_5117_32 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_5117_33 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_5117_34 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_5117_35 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_5117_36 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_5117_37 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_5117_38 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_5117_39 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_5117_40 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_5117_41 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_5117_42 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_5117_43 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_5117_44 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_5117_45 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_5117_46 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_5117_47 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_5117_48 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_5117_49 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_5117_50 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_5117_51 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_5117_52 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_5117_53 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_5117_54 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_5117_55 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_5117_56 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_5117_57 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_5117_58 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_5117_59 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_5117_60 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_5117_61 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_5117_62 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_5117_63 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_5581_0 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_5581_1 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_5581_2 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_5581_3 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_5581_4 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_5581_5 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_5581_6 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_5581_7 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_5581_8 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_5581_9 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_5581_10 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_5581_11 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_5581_12 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_5581_13 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_5581_14 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_5581_15 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_5581_16 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_5581_17 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_5581_18 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_5581_19 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_5581_20 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_5581_21 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_5581_22 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_5581_23 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_5581_24 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_5581_25 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_5581_26 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_5581_27 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_5581_28 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_5581_29 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_5581_30 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_5581_31 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_5581_32 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_5581_33 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_5581_34 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_5581_35 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_5581_36 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_5581_37 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_5581_38 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_5581_39 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_5581_40 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_5581_41 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_5581_42 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_5581_43 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_5581_44 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_5581_45 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_5581_46 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_5581_47 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_5581_48 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_5581_49 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_5581_50 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_5581_51 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_5581_52 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_5581_53 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_5581_54 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_5581_55 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_5581_56 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_5581_57 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_5581_58 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_5581_59 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_5581_60 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_5581_61 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_5581_62 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_5581_63 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5779 = _RAND_545[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5781 = _RAND_546[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5783 = _RAND_547[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5785 = _RAND_548[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5787 = _RAND_549[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_5789 = _RAND_550[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_5791 = _RAND_551[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_5793 = _RAND_552[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_5795 = _RAND_553[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_5797 = _RAND_554[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_5799 = _RAND_555[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_5801 = _RAND_556[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_5803 = _RAND_557[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_5805 = _RAND_558[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_5807 = _RAND_559[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_5809 = _RAND_560[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_5811 = _RAND_561[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_5813 = _RAND_562[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_5815 = _RAND_563[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_5817 = _RAND_564[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_5819 = _RAND_565[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_5821 = _RAND_566[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_5823 = _RAND_567[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_5825 = _RAND_568[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_5827 = _RAND_569[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_5829 = _RAND_570[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_5831 = _RAND_571[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_5833 = _RAND_572[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_5835 = _RAND_573[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_5837 = _RAND_574[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_5839 = _RAND_575[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_5841 = _RAND_576[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_5843 = _RAND_577[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_5845 = _RAND_578[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_5847 = _RAND_579[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_5849 = _RAND_580[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_5851 = _RAND_581[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_5853 = _RAND_582[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_5855 = _RAND_583[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_5857 = _RAND_584[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_5859 = _RAND_585[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_5861 = _RAND_586[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_5863 = _RAND_587[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_5865 = _RAND_588[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_5867 = _RAND_589[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_5869 = _RAND_590[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_5871 = _RAND_591[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_5873 = _RAND_592[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_5875 = _RAND_593[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_5877 = _RAND_594[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_5879 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_5881 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_5883 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_5885 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_5887 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_5889 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_5891 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_5893 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_5895 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_5897 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_5899 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_5901 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_5903 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_5905 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_5907 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_5909 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_5911 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_5913 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_5915 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_5917 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_5919 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_5921 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_5923 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_5925 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_5927 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_5929 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_5931 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_5933 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_5935 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_5937 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_5939 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_5941 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_5943 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_5945 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_5947 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_5949 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_5951 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_5953 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_5955 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_5957 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_5959 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_5961 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_5963 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_5965 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_5967 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_5969 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_5971 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_5973 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_5975 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_5977 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_5979 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_5981 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_5983 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_5985 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_5987 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_5989 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_5991 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_5993 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_5995 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_5997 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_5999 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_6001 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_6003 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_6005 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_6007 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_6009 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_6011 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_6013 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_6015 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_6017 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_6019 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_6021 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_6023 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_6025 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_6027 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_6029 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_6031 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_6033 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (_T_623) begin
      _T_718 <= 1'h0;
    end else begin
      _T_718 <= _T_633;
    end
    if (_T_623) begin
      _T_725 <= 6'h0;
    end else begin
      if (_T_633) begin
        _T_725 <= 6'h1;
      end
    end
    if (_T_623) begin
      _T_732 <= 14'h0;
    end else begin
      if (_T_633) begin
        _T_732 <= {{2'd0}, _T_808};
      end
    end
    if (_T_623) begin
      _T_739 <= 14'h0;
    end else begin
      if (_T_633) begin
        _T_739 <= {{2'd0}, _T_801};
      end
    end
    if (_T_623) begin
      _T_746 <= 15'h0;
    end else begin
      if (_T_633) begin
        _T_746 <= _T_797;
      end
    end
    if (_T_623) begin
      _T_753 <= 15'h0;
    end else begin
      if (_T_633) begin
        _T_753 <= _T_800;
      end
    end
    if (_T_623) begin
      _T_760 <= 13'h0;
    end else begin
      if (_T_633) begin
        _T_760 <= io_reg2dp_dataout_width;
      end
    end
    if (_T_623) begin
      _T_774 <= 15'h0;
    end else begin
      if (_T_718) begin
        _T_774 <= _T_816;
      end
    end
    if (_T_623) begin
      _T_781 <= 12'h0;
    end else begin
      if (_T_718) begin
        _T_781 <= _T_803;
      end
    end
    if (_T_623) begin
      _T_788 <= 12'h0;
    end else begin
      if (_T_718) begin
        _T_788 <= _T_805;
      end
    end
    if (_T_623) begin
      _T_795 <= 14'h0;
    end else begin
      if (_T_633) begin
        if (io_reg2dp_skip_data_rls) begin
          _T_795 <= _T_810;
        end else begin
          _T_795 <= _T_812;
        end
      end
    end
    if (_T_623) begin
      _T_834 <= 34'h0;
    end else begin
      if (_T_633) begin
        if (_T_638) begin
          _T_834 <= 34'h3ffffffff;
        end else begin
          _T_834 <= 34'h0;
        end
      end
    end
    if (_T_623) begin
      _T_841 <= 5'h0;
    end else begin
      if (_T_633) begin
        _T_841 <= _T_1044;
      end
    end
    if (_T_623) begin
      _T_848 <= 14'h0;
    end else begin
      if (_T_633) begin
        _T_848 <= _T_1046;
      end
    end
    if (_T_623) begin
      _T_855 <= 13'h0;
    end else begin
      if (_T_633) begin
        _T_855 <= io_reg2dp_datain_width_ext;
      end
    end
    if (_T_623) begin
      _T_862 <= 13'h0;
    end else begin
      if (_T_633) begin
        _T_862 <= io_reg2dp_datain_height_ext;
      end
    end
    if (_T_623) begin
      _T_869 <= 11'h0;
    end else begin
      if (_T_633) begin
        _T_869 <= _T_1053;
      end
    end
    if (_T_623) begin
      _T_872 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_872 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_875 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_875 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_881 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_881 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_884 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_884 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_887 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_887 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_890 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_890 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_896 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_896 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_899 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_899 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_905 <= 3'h1;
    end else begin
      if (_T_633) begin
        _T_905 <= _T_646;
      end
    end
    if (_T_623) begin
      _T_908 <= 3'h1;
    end else begin
      if (_T_633) begin
        if (_T_638) begin
          _T_908 <= _T_646;
        end else begin
          _T_908 <= 3'h1;
        end
      end
    end
    if (_T_623) begin
      _T_911 <= 3'h1;
    end else begin
      if (_T_633) begin
        if (_T_638) begin
          _T_911 <= _T_646;
        end else begin
          _T_911 <= 3'h1;
        end
      end
    end
    if (_T_623) begin
      _T_918 <= 4'h0;
    end else begin
      if (_T_633) begin
        _T_918 <= _T_653;
      end
    end
    if (_T_623) begin
      _T_925 <= 4'h0;
    end else begin
      if (_T_633) begin
        _T_925 <= _T_707;
      end
    end
    if (_T_623) begin
      _T_935 <= 5'h0;
    end else begin
      if (_T_633) begin
        _T_935 <= 5'h0;
      end
    end
    if (_T_623) begin
      _T_942 <= 7'h0;
    end else begin
      if (_T_633) begin
        if (_T_689) begin
          _T_942 <= _T_682;
        end else begin
          _T_942 <= {{1'd0}, _T_688};
        end
      end
    end
    if (_T_623) begin
      _T_949 <= 7'h0;
    end else begin
      if (_T_633) begin
        _T_949 <= _T_693;
      end
    end
    if (_T_623) begin
      _T_956 <= 8'h0;
    end else begin
      if (_T_633) begin
        if (_T_689) begin
          _T_956 <= _T_696;
        end else begin
          _T_956 <= {{1'd0}, _T_701};
        end
      end
    end
    if (_T_623) begin
      _T_963 <= 7'h0;
    end else begin
      if (_T_633) begin
        _T_963 <= {{1'd0}, _T_665};
      end
    end
    if (_T_623) begin
      _T_970 <= 12'h0;
    end else begin
      if (_T_633) begin
        _T_970 <= _T_705;
      end
    end
    if (_T_623) begin
      _T_977 <= 6'h0;
    end else begin
      if (_T_633) begin
        if (_T_638) begin
          _T_977 <= 6'h1;
        end else begin
          _T_977 <= _T_710;
        end
      end
    end
    if (_T_623) begin
      _T_984 <= 6'h0;
    end else begin
      if (_T_633) begin
        if (_T_638) begin
          _T_984 <= 6'h1;
        end else begin
          _T_984 <= _T_714;
        end
      end
    end
    if (_T_623) begin
      _T_991 <= 16'h0;
    end else begin
      if (_T_633) begin
        _T_991 <= io_reg2dp_pad_value;
      end
    end
    if (_T_623) begin
      _T_998 <= 15'h0;
    end else begin
      if (_T_633) begin
        _T_998 <= _T_1057;
      end
    end
    if (_T_623) begin
      _T_1005 <= 15'h0;
    end else begin
      if (_T_718) begin
        _T_1005 <= _T_746;
      end
    end
    if (_T_623) begin
      _T_1012 <= 15'h0;
    end else begin
      if (_T_718) begin
        _T_1012 <= _T_746;
      end
    end
    if (_T_623) begin
      _T_1019 <= 14'h0;
    end else begin
      if (_T_629) begin
        _T_1019 <= _T_795;
      end
    end
    if (_T_623) begin
      _T_1026 <= 15'h0;
    end else begin
      if (_T_629) begin
        _T_1026 <= _T_816;
      end
    end
    if (_T_623) begin
      _T_2220 <= 1'h0;
    end else begin
      _T_2220 <= _T_2217;
    end
    if (_T_623) begin
      _T_2214 <= 1'h0;
    end else begin
      _T_2214 <= _T_2211;
    end
    if (_T_623) begin
      _T_2211 <= 1'h0;
    end else begin
      _T_2211 <= _T_1961;
    end
    if (_T_623) begin
      _T_2234 <= 27'h0;
    end else begin
      if (_T_2217) begin
        _T_2234 <= _T_2231;
      end
    end
    if (_T_623) begin
      _T_2228 <= 27'h0;
    end else begin
      if (_T_2211) begin
        _T_2228 <= _T_2225;
      end
    end
    if (_T_623) begin
      _T_2225 <= 27'h0;
    end else begin
      if (_T_1961) begin
        _T_2225 <= _T_2243;
      end
    end
    if (_T_623) begin
      _T_1169 <= 1'h0;
    end else begin
      _T_1169 <= _T_1164;
    end
    if (_T_623) begin
      _T_1172 <= 14'h0;
    end else begin
      if (_T_1164) begin
        if (_T_1157) begin
          _T_1172 <= _T_732;
        end else begin
          _T_1172 <= _T_1019;
        end
      end
    end
    if (_T_623) begin
      _T_1175 <= 15'h0;
    end else begin
      if (_T_1164) begin
        if (_T_1157) begin
          _T_1175 <= _T_774;
        end else begin
          _T_1175 <= _T_1026;
        end
      end
    end
    if (_T_623) begin
      _T_1180 <= 1'h0;
    end else begin
      _T_1180 <= io_sg2dl_pd_valid;
    end
    if (_T_623) begin
      _T_1183 <= 1'h0;
    end else begin
      _T_1183 <= _T_1180;
    end
    if (_T_623) begin
      _T_1186 <= 1'h0;
    end else begin
      _T_1186 <= _T_1183;
    end
    if (_T_623) begin
      _T_1189 <= 1'h0;
    end else begin
      _T_1189 <= _T_1186;
    end
    if (_T_623) begin
      _T_1192 <= 1'h0;
    end else begin
      _T_1192 <= _T_1189;
    end
    if (_T_623) begin
      _T_1214 <= 1'h0;
    end else begin
      _T_1214 <= _T_1192;
    end
    if (_T_623) begin
      _T_1217 <= 1'h0;
    end else begin
      _T_1217 <= _T_1214;
    end
    if (_T_623) begin
      _T_1220 <= 1'h0;
    end else begin
      _T_1220 <= _T_1217;
    end
    if (_T_623) begin
      _T_1223 <= 1'h0;
    end else begin
      _T_1223 <= _T_1220;
    end
    if (_T_623) begin
      _T_1228 <= 31'h0;
    end else begin
      if (_T_1192) begin
        _T_1228 <= _T_1225;
      end
    end
    if (_T_623) begin
      _T_1231 <= 31'h0;
    end else begin
      if (_T_1214) begin
        _T_1231 <= _T_1228;
      end
    end
    if (_T_623) begin
      _T_1234 <= 31'h0;
    end else begin
      if (_T_1217) begin
        _T_1234 <= _T_1231;
      end
    end
    if (_T_623) begin
      _T_1237 <= 31'h0;
    end else begin
      if (_T_1220) begin
        _T_1237 <= _T_1234;
      end
    end
    if (_T_623) begin
      _T_1282 <= 5'h0;
    end else begin
      if (_T_633) begin
        _T_1282 <= 5'h0;
      end else begin
        if (_T_1290) begin
          _T_1282 <= 5'h0;
        end else begin
          _T_1282 <= _T_1287;
        end
      end
    end
    if (_T_623) begin
      _T_1293 <= 2'h0;
    end else begin
      if (_T_1303) begin
        if (_T_1304) begin
          _T_1293 <= 2'h0;
        end else begin
          _T_1293 <= _T_1298;
        end
      end
    end
    if (_T_623) begin
      _T_1309 <= 7'h0;
    end else begin
      if (_T_1321) begin
        if (_T_633) begin
          _T_1309 <= 7'h0;
        end else begin
          if (_T_1324) begin
            _T_1309 <= 7'h0;
          end else begin
            if (_T_1319) begin
              _T_1309 <= 7'h0;
            end else begin
              _T_1309 <= _T_1316;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1338 <= 1'h0;
    end else begin
      if (_T_1245) begin
        _T_1338 <= 1'h1;
      end else begin
        if (_T_1358) begin
          _T_1338 <= 1'h0;
        end
      end
    end
    if (_T_623) begin
      _T_1332 <= 1'h0;
    end else begin
      if (_T_1341) begin
        _T_1332 <= 1'h0;
      end else begin
        if (_T_1245) begin
          _T_1332 <= 1'h1;
        end
      end
    end
    if (_T_623) begin
      _T_1335 <= 1'h0;
    end else begin
      _T_1335 <= _T_1346;
    end
    if (_T_623) begin
      _T_1364 <= 8'h0;
    end else begin
      if (_T_1361) begin
        _T_1364 <= _T_1366;
      end
    end
    if (_T_623) begin
      _T_1369 <= 13'h0;
    end else begin
      if (_T_1387) begin
        if (_T_633) begin
          _T_1369 <= {{9'd0}, _T_651};
        end else begin
          if (_T_1381) begin
            _T_1369 <= _T_1372;
          end else begin
            if (_T_1377) begin
              _T_1369 <= {{9'd0}, _T_651};
            end else begin
              _T_1369 <= _T_1374;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1372 <= 13'h0;
    end else begin
      if (_T_1390) begin
        if (_T_633) begin
          _T_1372 <= {{9'd0}, _T_651};
        end else begin
          if (!(_T_1381)) begin
            if (_T_1377) begin
              _T_1372 <= {{9'd0}, _T_651};
            end else begin
              _T_1372 <= _T_1374;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1393 <= 11'h0;
    end else begin
      if (_T_1397) begin
        if (_T_633) begin
          _T_1393 <= 11'h0;
        end else begin
          if (_T_1272) begin
            _T_1393 <= 11'h0;
          end else begin
            _T_1393 <= _T_1402;
          end
        end
      end
    end
    if (_T_623) begin
      _T_1407 <= 14'h0;
    end else begin
      if (_T_1451) begin
        if (_T_633) begin
          if (_T_638) begin
            _T_1407 <= 14'h0;
          end else begin
            _T_1407 <= _T_1434;
          end
        end else begin
          if (_T_1381) begin
            _T_1407 <= _T_1410;
          end else begin
            if (_T_1377) begin
              if (_T_638) begin
                _T_1407 <= 14'h0;
              end else begin
                _T_1407 <= _T_1434;
              end
            end else begin
              _T_1407 <= _T_1437;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1410 <= 14'h0;
    end else begin
      if (_T_1457) begin
        if (_T_633) begin
          if (_T_638) begin
            _T_1410 <= 14'h0;
          end else begin
            _T_1410 <= _T_1434;
          end
        end else begin
          if (!(_T_1381)) begin
            if (_T_1377) begin
              if (_T_638) begin
                _T_1410 <= 14'h0;
              end else begin
                _T_1410 <= _T_1434;
              end
            end else begin
              _T_1410 <= _T_1437;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1413 <= 16'h0;
    end else begin
      if (_T_1451) begin
        if (_T_718) begin
          _T_1413 <= {{9'd0}, _T_942};
        end else begin
          if (_T_1480) begin
            _T_1413 <= {{9'd0}, _T_942};
          end else begin
            if (_T_1484) begin
              _T_1413 <= _T_1486;
            end else begin
              if (_T_1488) begin
                _T_1413 <= _T_1490;
              end else begin
                if (_T_1493) begin
                  _T_1413 <= _T_1496;
                end else begin
                  if (_T_1498) begin
                    _T_1413 <= _T_1416;
                  end else begin
                    _T_1413 <= _T_1500;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1416 <= 16'h0;
    end else begin
      if (_T_1457) begin
        if (_T_718) begin
          _T_1416 <= {{9'd0}, _T_942};
        end else begin
          if (_T_1480) begin
            _T_1416 <= {{9'd0}, _T_942};
          end else begin
            if (_T_1484) begin
              _T_1416 <= _T_1486;
            end else begin
              if (_T_1488) begin
                _T_1416 <= _T_1490;
              end else begin
                if (_T_1493) begin
                  _T_1416 <= _T_1496;
                end else begin
                  if (!(_T_1498)) begin
                    _T_1416 <= _T_1500;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1419 <= 16'h0;
    end else begin
      if (_T_1529) begin
        if (_T_718) begin
          _T_1419 <= {{9'd0}, _T_942};
        end else begin
          if (_T_1480) begin
            _T_1419 <= {{9'd0}, _T_942};
          end else begin
            if (_T_1484) begin
              _T_1419 <= _T_1486;
            end else begin
              if (_T_1488) begin
                _T_1419 <= _T_1490;
              end else begin
                if (_T_1493) begin
                  _T_1419 <= _T_1496;
                end else begin
                  if (_T_1498) begin
                    _T_1419 <= _T_1416;
                  end else begin
                    _T_1419 <= _T_1500;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1422 <= 13'h2;
    end else begin
      if (_T_1469) begin
        _T_1422 <= 13'h2;
      end else begin
        if (_T_1471) begin
          _T_1422 <= _T_1474;
        end
      end
    end
    if (_T_623) begin
      _T_1427 <= 1'h0;
    end else begin
      if (_T_1361) begin
        _T_1427 <= _T_1539;
      end
    end
    if (_T_623) begin
      _T_1430 <= 1'h0;
    end else begin
      if (_T_1361) begin
        if (_T_1531) begin
          _T_1430 <= 1'h1;
        end else begin
          if (_T_1427) begin
            _T_1430 <= 1'h0;
          end
        end
      end
    end
    if (_T_623) begin
      _T_1542 <= 14'h0;
    end else begin
      if (_T_1563) begin
        if (_T_1553) begin
          _T_1542 <= _T_1549;
        end else begin
          if (_T_1381) begin
            _T_1542 <= _T_1545;
          end else begin
            if (_T_1377) begin
              _T_1542 <= _T_1551;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1545 <= 14'h0;
    end else begin
      if (_T_1390) begin
        if (_T_1553) begin
          _T_1545 <= _T_1549;
        end else begin
          if (!(_T_1381)) begin
            if (_T_1377) begin
              _T_1545 <= _T_1551;
            end else begin
              _T_1545 <= _T_1542;
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_1619 <= 1'h0;
    end else begin
      _T_1619 <= _T_1603;
    end
    if (_T_623) begin
      _T_1622 <= 2'h0;
    end else begin
      if (_T_1361) begin
        _T_1622 <= _T_1608;
      end
    end
    if (_T_623) begin
      _T_1625 <= 2'h0;
    end else begin
      if (_T_1361) begin
        _T_1625 <= _T_1293;
      end
    end
    if (_T_623) begin
      _T_1628 <= 1'h0;
    end else begin
      if (_T_1361) begin
        if (_T_1605) begin
          _T_1628 <= _T_1606;
        end else begin
          _T_1628 <= _T_1271;
        end
      end
    end
    if (_T_623) begin
      _T_1631 <= 1'h0;
    end else begin
      if (_T_1361) begin
        _T_1631 <= _T_1394;
      end
    end
    if (_T_623) begin
      _T_1634 <= 1'h0;
    end else begin
      if (_T_1361) begin
        if (_T_1245) begin
          _T_1634 <= 1'h1;
        end else begin
          if (_T_1358) begin
            _T_1634 <= 1'h0;
          end else begin
            _T_1634 <= _T_1338;
          end
        end
      end
    end
    if (_T_623) begin
      _T_1637 <= 2'h0;
    end else begin
      if (_T_1361) begin
        _T_1637 <= _T_1270;
      end
    end
    if (_T_623) begin
      _T_1640 <= 1'h0;
    end else begin
      if (_T_1611) begin
        _T_1640 <= _T_1245;
      end
    end
    if (_T_623) begin
      _T_1643 <= 9'h0;
    end else begin
      if (_T_1361) begin
        _T_1643 <= _T_1616;
      end
    end
    if (_T_623) begin
      _T_1646 <= 1'h0;
    end else begin
      if (_T_1361) begin
        _T_1646 <= _T_1648;
      end
    end
    if (_T_623) begin
      _T_1651 <= 13'h0;
    end else begin
      if (_T_1397) begin
        if (_T_633) begin
          _T_1651 <= 13'h0;
        end else begin
          if (_T_1676) begin
            _T_1651 <= 13'h0;
          end else begin
            _T_1651 <= _T_1679;
          end
        end
      end
    end
    if (_T_623) begin
      _T_1654 <= 13'h0;
    end else begin
      if (_T_1685) begin
        _T_1654 <= _T_1651;
      end
    end
    if (_T_623) begin
      _T_1657 <= 13'h0;
    end else begin
      if (_T_1718) begin
        _T_1657 <= _T_1687;
      end
    end
    if (_T_623) begin
      _T_1660 <= 13'h0;
    end else begin
      if (_T_1718) begin
        _T_1660 <= _T_1689;
      end
    end
    if (_T_623) begin
      _T_1663 <= 13'h0;
    end else begin
      if (_T_1718) begin
        _T_1663 <= _T_1691;
      end
    end
    if (_T_623) begin
      _T_1666 <= 13'h0;
    end else begin
      if (_T_1719) begin
        _T_1666 <= _T_1695;
      end
    end
    if (_T_623) begin
      _T_1669 <= 13'h0;
    end else begin
      _T_1669 <= _GEN_95[12:0];
    end
    if (_T_623) begin
      _T_1762_0 <= 13'h1fff;
    end else begin
      _T_1762_0 <= _GEN_96[12:0];
    end
    if (_T_623) begin
      _T_1762_1 <= 13'h1fff;
    end else begin
      _T_1762_1 <= _GEN_97[12:0];
    end
    if (_T_623) begin
      _T_1762_2 <= 13'h1fff;
    end else begin
      _T_1762_2 <= _GEN_98[12:0];
    end
    if (_T_623) begin
      _T_1762_3 <= 13'h1fff;
    end else begin
      _T_1762_3 <= _GEN_99[12:0];
    end
    if (_T_623) begin
      _T_1781 <= 1'h0;
    end else begin
      _T_1781 <= _T_1894;
    end
    if (_T_623) begin
      _T_1788 <= 15'h1fff;
    end else begin
      if (_T_1925) begin
        if (_T_1853) begin
          _T_1788 <= 15'h1fff;
        end else begin
          if (_T_1843) begin
            _T_1788 <= _T_1852;
          end else begin
            _T_1788 <= _T_1836;
          end
        end
      end
    end
    if (_T_623) begin
      _T_1791 <= 1'h0;
    end else begin
      _T_1791 <= _T_1335;
    end
    if (_T_623) begin
      _T_1797 <= 2'h0;
    end else begin
      if (_T_1338) begin
        _T_1797 <= _T_1622;
      end
    end
    if (_T_623) begin
      _T_1800 <= 2'h0;
    end else begin
      if (_T_1338) begin
        _T_1800 <= _T_1625;
      end
    end
    if (_T_623) begin
      _T_1803 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1803 <= _T_1628;
      end
    end
    if (_T_623) begin
      _T_1806 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1806 <= _T_1631;
      end
    end
    if (_T_623) begin
      _T_1809 <= 8'h0;
    end else begin
      if (_T_1338) begin
        _T_1809 <= _T_1364;
      end
    end
    if (_T_623) begin
      _T_1812 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1812 <= _T_1634;
      end
    end
    if (_T_623) begin
      _T_1815 <= 2'h0;
    end else begin
      if (_T_1338) begin
        _T_1815 <= _T_1637;
      end
    end
    if (_T_623) begin
      _T_1818 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1818 <= _T_1640;
      end
    end
    if (_T_623) begin
      _T_1821 <= 1'h0;
    end else begin
      if (_T_1338) begin
        _T_1821 <= _T_1646;
      end
    end
    if (_T_623) begin
      _T_1824 <= 9'h0;
    end else begin
      if (_T_1338) begin
        _T_1824 <= _T_1643;
      end else begin
        _T_1824 <= {{8'd0}, _T_1338};
      end
    end
    if (_T_623) begin
      _T_1946 <= 1'h0;
    end else begin
      _T_1946 <= _T_1791;
    end
    if (_T_623) begin
      _T_1949 <= 1'h0;
    end else begin
      _T_1949 <= _T_1946;
    end
    if (_T_623) begin
      _T_1952 <= 1'h0;
    end else begin
      _T_1952 <= _T_1949;
    end
    if (_T_623) begin
      _T_1955 <= 1'h0;
    end else begin
      _T_1955 <= _T_1952;
    end
    if (_T_623) begin
      _T_1958 <= 1'h0;
    end else begin
      _T_1958 <= _T_1955;
    end
    if (_T_623) begin
      _T_1961 <= 1'h0;
    end else begin
      _T_1961 <= _T_1958;
    end
    if (_T_623) begin
      _T_1966 <= 29'h0;
    end else begin
      if (_T_1791) begin
        _T_1966 <= _T_1941;
      end
    end
    if (_T_623) begin
      _T_1969 <= 29'h0;
    end else begin
      if (_T_1946) begin
        _T_1969 <= _T_1966;
      end
    end
    if (_T_623) begin
      _T_1972 <= 29'h0;
    end else begin
      if (_T_1949) begin
        _T_1972 <= _T_1969;
      end
    end
    if (_T_623) begin
      _T_1975 <= 29'h0;
    end else begin
      if (_T_1952) begin
        _T_1975 <= _T_1972;
      end
    end
    if (_T_623) begin
      _T_1978 <= 29'h0;
    end else begin
      if (_T_1955) begin
        _T_1978 <= _T_1975;
      end
    end
    if (_T_623) begin
      _T_1981 <= 29'h0;
    end else begin
      if (_T_1958) begin
        _T_1981 <= _T_1978;
      end
    end
    if (_T_623) begin
      _T_2054 <= 1'h1;
    end else begin
      if (io_sc2buf_dat_rd_data_valid) begin
        _T_2054 <= 1'h0;
      end
    end
    if (_T_623) begin
      _T_2066 <= 1'h1;
    end else begin
      if (_T_2111) begin
        _T_2066 <= 1'h0;
      end else begin
        if (io_sc2buf_dat_rd_data_valid) begin
          _T_2066 <= _T_2054;
        end
      end
    end
    if (io_sc2buf_dat_rd_data_valid) begin
      _T_2077 <= io_sc2buf_dat_rd_data_bits;
    end
    if (_T_2111) begin
      _T_2085 <= _T_2077;
    end
    if (_T_623) begin
      _T_2185 <= 8'h0;
    end else begin
      if (_T_2391) begin
        if (_T_633) begin
          _T_2185 <= 8'h40;
        end else begin
          if (_T_2347) begin
            _T_2185 <= _T_2197;
          end else begin
            if (_T_2348) begin
              _T_2185 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2185 <= 8'h40;
              end else begin
                _T_2185 <= _T_2316;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2188 <= 8'h0;
    end else begin
      if (_T_2397) begin
        if (_T_633) begin
          _T_2188 <= 8'h40;
        end else begin
          if (_T_2358) begin
            _T_2188 <= _T_2200;
          end else begin
            if (_T_2359) begin
              _T_2188 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2188 <= 8'h40;
              end else begin
                _T_2188 <= _T_2325;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2191 <= 8'h0;
    end else begin
      if (_T_2403) begin
        if (_T_633) begin
          _T_2191 <= 8'h40;
        end else begin
          if (_T_2369) begin
            _T_2191 <= _T_2203;
          end else begin
            if (_T_2370) begin
              _T_2191 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2191 <= 8'h40;
              end else begin
                _T_2191 <= _T_2334;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2194 <= 8'h0;
    end else begin
      if (_T_2409) begin
        if (_T_633) begin
          _T_2194 <= 8'h40;
        end else begin
          if (_T_2380) begin
            _T_2194 <= _T_2206;
          end else begin
            if (_T_2381) begin
              _T_2194 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2194 <= 8'h40;
              end else begin
                _T_2194 <= _T_2343;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2197 <= 8'h0;
    end else begin
      if (_T_2414) begin
        if (_T_633) begin
          _T_2197 <= 8'h40;
        end else begin
          if (!(_T_2347)) begin
            if (_T_2348) begin
              _T_2197 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2197 <= 8'h40;
              end else begin
                _T_2197 <= _T_2316;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2200 <= 8'h0;
    end else begin
      if (_T_2422) begin
        if (_T_633) begin
          _T_2200 <= 8'h40;
        end else begin
          if (!(_T_2358)) begin
            if (_T_2359) begin
              _T_2200 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2200 <= 8'h40;
              end else begin
                _T_2200 <= _T_2325;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2203 <= 8'h0;
    end else begin
      if (_T_2430) begin
        if (_T_633) begin
          _T_2203 <= 8'h40;
        end else begin
          if (!(_T_2369)) begin
            if (_T_2370) begin
              _T_2203 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2203 <= 8'h40;
              end else begin
                _T_2203 <= _T_2334;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2206 <= 8'h0;
    end else begin
      if (_T_2438) begin
        if (_T_633) begin
          _T_2206 <= 8'h40;
        end else begin
          if (!(_T_2380)) begin
            if (_T_2381) begin
              _T_2206 <= 8'h40;
            end else begin
              if (_T_2310) begin
                _T_2206 <= 8'h40;
              end else begin
                _T_2206 <= _T_2343;
              end
            end
          end
        end
      end
    end
    if (_T_623) begin
      _T_2217 <= 1'h0;
    end else begin
      _T_2217 <= _T_2214;
    end
    if (_T_623) begin
      _T_2231 <= 27'h0;
    end else begin
      if (_T_2214) begin
        _T_2231 <= _T_2228;
      end
    end
    _T_2614 <= _GEN_149[255:0];
    _T_2616 <= _GEN_150[127:0];
    if (_T_2824) begin
      _T_2618 <= _T_2616;
    end
    _T_2620 <= _GEN_151[127:0];
    if (_T_2824) begin
      _T_2622 <= _T_2620;
    end
    _T_2624 <= _GEN_154[127:0];
    if (_T_623) begin
      _T_3422 <= 1'h0;
    end else begin
      _T_3422 <= _T_2251;
    end
    if (_T_623) begin
      _T_3692_0 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_0 <= _T_3223;
      end
    end
    if (_T_623) begin
      _T_3692_1 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_1 <= _T_3225;
      end
    end
    if (_T_623) begin
      _T_3692_2 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_2 <= _T_3227;
      end
    end
    if (_T_623) begin
      _T_3692_3 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_3 <= _T_3229;
      end
    end
    if (_T_623) begin
      _T_3692_4 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_4 <= _T_3231;
      end
    end
    if (_T_623) begin
      _T_3692_5 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_5 <= _T_3233;
      end
    end
    if (_T_623) begin
      _T_3692_6 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_6 <= _T_3235;
      end
    end
    if (_T_623) begin
      _T_3692_7 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_7 <= _T_3237;
      end
    end
    if (_T_623) begin
      _T_3692_8 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_8 <= _T_3239;
      end
    end
    if (_T_623) begin
      _T_3692_9 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_9 <= _T_3241;
      end
    end
    if (_T_623) begin
      _T_3692_10 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_10 <= _T_3243;
      end
    end
    if (_T_623) begin
      _T_3692_11 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_11 <= _T_3245;
      end
    end
    if (_T_623) begin
      _T_3692_12 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_12 <= _T_3247;
      end
    end
    if (_T_623) begin
      _T_3692_13 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_13 <= _T_3249;
      end
    end
    if (_T_623) begin
      _T_3692_14 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_14 <= _T_3251;
      end
    end
    if (_T_623) begin
      _T_3692_15 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_15 <= _T_3253;
      end
    end
    if (_T_623) begin
      _T_3692_16 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_16 <= _T_3255;
      end
    end
    if (_T_623) begin
      _T_3692_17 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_17 <= _T_3257;
      end
    end
    if (_T_623) begin
      _T_3692_18 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_18 <= _T_3259;
      end
    end
    if (_T_623) begin
      _T_3692_19 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_19 <= _T_3261;
      end
    end
    if (_T_623) begin
      _T_3692_20 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_20 <= _T_3263;
      end
    end
    if (_T_623) begin
      _T_3692_21 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_21 <= _T_3265;
      end
    end
    if (_T_623) begin
      _T_3692_22 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_22 <= _T_3267;
      end
    end
    if (_T_623) begin
      _T_3692_23 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_23 <= _T_3269;
      end
    end
    if (_T_623) begin
      _T_3692_24 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_24 <= _T_3271;
      end
    end
    if (_T_623) begin
      _T_3692_25 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_25 <= _T_3273;
      end
    end
    if (_T_623) begin
      _T_3692_26 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_26 <= _T_3275;
      end
    end
    if (_T_623) begin
      _T_3692_27 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_27 <= _T_3277;
      end
    end
    if (_T_623) begin
      _T_3692_28 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_28 <= _T_3279;
      end
    end
    if (_T_623) begin
      _T_3692_29 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_29 <= _T_3281;
      end
    end
    if (_T_623) begin
      _T_3692_30 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_30 <= _T_3283;
      end
    end
    if (_T_623) begin
      _T_3692_31 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_31 <= _T_3285;
      end
    end
    if (_T_623) begin
      _T_3692_32 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_32 <= _T_3287;
      end
    end
    if (_T_623) begin
      _T_3692_33 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_33 <= _T_3289;
      end
    end
    if (_T_623) begin
      _T_3692_34 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_34 <= _T_3291;
      end
    end
    if (_T_623) begin
      _T_3692_35 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_35 <= _T_3293;
      end
    end
    if (_T_623) begin
      _T_3692_36 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_36 <= _T_3295;
      end
    end
    if (_T_623) begin
      _T_3692_37 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_37 <= _T_3297;
      end
    end
    if (_T_623) begin
      _T_3692_38 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_38 <= _T_3299;
      end
    end
    if (_T_623) begin
      _T_3692_39 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_39 <= _T_3301;
      end
    end
    if (_T_623) begin
      _T_3692_40 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_40 <= _T_3303;
      end
    end
    if (_T_623) begin
      _T_3692_41 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_41 <= _T_3305;
      end
    end
    if (_T_623) begin
      _T_3692_42 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_42 <= _T_3307;
      end
    end
    if (_T_623) begin
      _T_3692_43 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_43 <= _T_3309;
      end
    end
    if (_T_623) begin
      _T_3692_44 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_44 <= _T_3311;
      end
    end
    if (_T_623) begin
      _T_3692_45 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_45 <= _T_3313;
      end
    end
    if (_T_623) begin
      _T_3692_46 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_46 <= _T_3315;
      end
    end
    if (_T_623) begin
      _T_3692_47 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_47 <= _T_3317;
      end
    end
    if (_T_623) begin
      _T_3692_48 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_48 <= _T_3319;
      end
    end
    if (_T_623) begin
      _T_3692_49 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_49 <= _T_3321;
      end
    end
    if (_T_623) begin
      _T_3692_50 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_50 <= _T_3323;
      end
    end
    if (_T_623) begin
      _T_3692_51 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_51 <= _T_3325;
      end
    end
    if (_T_623) begin
      _T_3692_52 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_52 <= _T_3327;
      end
    end
    if (_T_623) begin
      _T_3692_53 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_53 <= _T_3329;
      end
    end
    if (_T_623) begin
      _T_3692_54 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_54 <= _T_3331;
      end
    end
    if (_T_623) begin
      _T_3692_55 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_55 <= _T_3333;
      end
    end
    if (_T_623) begin
      _T_3692_56 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_56 <= _T_3335;
      end
    end
    if (_T_623) begin
      _T_3692_57 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_57 <= _T_3337;
      end
    end
    if (_T_623) begin
      _T_3692_58 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_58 <= _T_3339;
      end
    end
    if (_T_623) begin
      _T_3692_59 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_59 <= _T_3341;
      end
    end
    if (_T_623) begin
      _T_3692_60 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_60 <= _T_3343;
      end
    end
    if (_T_623) begin
      _T_3692_61 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_61 <= _T_3345;
      end
    end
    if (_T_623) begin
      _T_3692_62 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_62 <= _T_3347;
      end
    end
    if (_T_623) begin
      _T_3692_63 <= 1'h0;
    end else begin
      if (_T_2251) begin
        _T_3692_63 <= _T_3349;
      end
    end
    if (_T_3959) begin
      if (_T_2891) begin
        _T_3892_0 <= _T_2752;
      end else begin
        _T_3892_0 <= _T_2549;
      end
    end
    if (_T_3960) begin
      if (_T_2891) begin
        _T_3892_1 <= _T_2753;
      end else begin
        _T_3892_1 <= _T_2550;
      end
    end
    if (_T_3961) begin
      if (_T_2891) begin
        _T_3892_2 <= _T_2754;
      end else begin
        _T_3892_2 <= _T_2551;
      end
    end
    if (_T_3962) begin
      if (_T_2891) begin
        _T_3892_3 <= _T_2755;
      end else begin
        _T_3892_3 <= _T_2552;
      end
    end
    if (_T_3963) begin
      if (_T_2891) begin
        _T_3892_4 <= _T_2756;
      end else begin
        _T_3892_4 <= _T_2553;
      end
    end
    if (_T_3964) begin
      if (_T_2891) begin
        _T_3892_5 <= _T_2757;
      end else begin
        _T_3892_5 <= _T_2554;
      end
    end
    if (_T_3965) begin
      if (_T_2891) begin
        _T_3892_6 <= _T_2758;
      end else begin
        _T_3892_6 <= _T_2555;
      end
    end
    if (_T_3966) begin
      if (_T_2891) begin
        _T_3892_7 <= _T_2759;
      end else begin
        _T_3892_7 <= _T_2556;
      end
    end
    if (_T_3967) begin
      if (_T_2891) begin
        _T_3892_8 <= _T_2760;
      end else begin
        _T_3892_8 <= _T_2557;
      end
    end
    if (_T_3968) begin
      if (_T_2891) begin
        _T_3892_9 <= _T_2761;
      end else begin
        _T_3892_9 <= _T_2558;
      end
    end
    if (_T_3969) begin
      if (_T_2891) begin
        _T_3892_10 <= _T_2762;
      end else begin
        _T_3892_10 <= _T_2559;
      end
    end
    if (_T_3970) begin
      if (_T_2891) begin
        _T_3892_11 <= _T_2763;
      end else begin
        _T_3892_11 <= _T_2560;
      end
    end
    if (_T_3971) begin
      if (_T_2891) begin
        _T_3892_12 <= _T_2764;
      end else begin
        _T_3892_12 <= _T_2561;
      end
    end
    if (_T_3972) begin
      if (_T_2891) begin
        _T_3892_13 <= _T_2765;
      end else begin
        _T_3892_13 <= _T_2562;
      end
    end
    if (_T_3973) begin
      if (_T_2891) begin
        _T_3892_14 <= _T_2766;
      end else begin
        _T_3892_14 <= _T_2563;
      end
    end
    if (_T_3974) begin
      if (_T_2891) begin
        _T_3892_15 <= _T_2767;
      end else begin
        _T_3892_15 <= _T_2564;
      end
    end
    if (_T_3975) begin
      if (_T_2891) begin
        _T_3892_16 <= _T_2768;
      end else begin
        _T_3892_16 <= _T_2565;
      end
    end
    if (_T_3976) begin
      if (_T_2891) begin
        _T_3892_17 <= _T_2769;
      end else begin
        _T_3892_17 <= _T_2566;
      end
    end
    if (_T_3977) begin
      if (_T_2891) begin
        _T_3892_18 <= _T_2770;
      end else begin
        _T_3892_18 <= _T_2567;
      end
    end
    if (_T_3978) begin
      if (_T_2891) begin
        _T_3892_19 <= _T_2771;
      end else begin
        _T_3892_19 <= _T_2568;
      end
    end
    if (_T_3979) begin
      if (_T_2891) begin
        _T_3892_20 <= _T_2772;
      end else begin
        _T_3892_20 <= _T_2569;
      end
    end
    if (_T_3980) begin
      if (_T_2891) begin
        _T_3892_21 <= _T_2773;
      end else begin
        _T_3892_21 <= _T_2570;
      end
    end
    if (_T_3981) begin
      if (_T_2891) begin
        _T_3892_22 <= _T_2774;
      end else begin
        _T_3892_22 <= _T_2571;
      end
    end
    if (_T_3982) begin
      if (_T_2891) begin
        _T_3892_23 <= _T_2775;
      end else begin
        _T_3892_23 <= _T_2572;
      end
    end
    if (_T_3983) begin
      if (_T_2891) begin
        _T_3892_24 <= _T_2776;
      end else begin
        _T_3892_24 <= _T_2573;
      end
    end
    if (_T_3984) begin
      if (_T_2891) begin
        _T_3892_25 <= _T_2777;
      end else begin
        _T_3892_25 <= _T_2574;
      end
    end
    if (_T_3985) begin
      if (_T_2891) begin
        _T_3892_26 <= _T_2778;
      end else begin
        _T_3892_26 <= _T_2575;
      end
    end
    if (_T_3986) begin
      if (_T_2891) begin
        _T_3892_27 <= _T_2779;
      end else begin
        _T_3892_27 <= _T_2576;
      end
    end
    if (_T_3987) begin
      if (_T_2891) begin
        _T_3892_28 <= _T_2780;
      end else begin
        _T_3892_28 <= _T_2577;
      end
    end
    if (_T_3988) begin
      if (_T_2891) begin
        _T_3892_29 <= _T_2781;
      end else begin
        _T_3892_29 <= _T_2578;
      end
    end
    if (_T_3989) begin
      if (_T_2891) begin
        _T_3892_30 <= _T_2782;
      end else begin
        _T_3892_30 <= _T_2579;
      end
    end
    if (_T_3990) begin
      if (_T_2891) begin
        _T_3892_31 <= _T_2783;
      end else begin
        _T_3892_31 <= _T_2580;
      end
    end
    if (_T_3991) begin
      if (_T_2891) begin
        _T_3892_32 <= _T_2784;
      end else begin
        _T_3892_32 <= _T_2581;
      end
    end
    if (_T_3992) begin
      if (_T_2891) begin
        _T_3892_33 <= _T_2785;
      end else begin
        _T_3892_33 <= _T_2582;
      end
    end
    if (_T_3993) begin
      if (_T_2891) begin
        _T_3892_34 <= _T_2786;
      end else begin
        _T_3892_34 <= _T_2583;
      end
    end
    if (_T_3994) begin
      if (_T_2891) begin
        _T_3892_35 <= _T_2787;
      end else begin
        _T_3892_35 <= _T_2584;
      end
    end
    if (_T_3995) begin
      if (_T_2891) begin
        _T_3892_36 <= _T_2788;
      end else begin
        _T_3892_36 <= _T_2585;
      end
    end
    if (_T_3996) begin
      if (_T_2891) begin
        _T_3892_37 <= _T_2789;
      end else begin
        _T_3892_37 <= _T_2586;
      end
    end
    if (_T_3997) begin
      if (_T_2891) begin
        _T_3892_38 <= _T_2790;
      end else begin
        _T_3892_38 <= _T_2587;
      end
    end
    if (_T_3998) begin
      if (_T_2891) begin
        _T_3892_39 <= _T_2791;
      end else begin
        _T_3892_39 <= _T_2588;
      end
    end
    if (_T_3999) begin
      if (_T_2891) begin
        _T_3892_40 <= _T_2792;
      end else begin
        _T_3892_40 <= _T_2589;
      end
    end
    if (_T_4000) begin
      if (_T_2891) begin
        _T_3892_41 <= _T_2793;
      end else begin
        _T_3892_41 <= _T_2590;
      end
    end
    if (_T_4001) begin
      if (_T_2891) begin
        _T_3892_42 <= _T_2794;
      end else begin
        _T_3892_42 <= _T_2591;
      end
    end
    if (_T_4002) begin
      if (_T_2891) begin
        _T_3892_43 <= _T_2795;
      end else begin
        _T_3892_43 <= _T_2592;
      end
    end
    if (_T_4003) begin
      if (_T_2891) begin
        _T_3892_44 <= _T_2796;
      end else begin
        _T_3892_44 <= _T_2593;
      end
    end
    if (_T_4004) begin
      if (_T_2891) begin
        _T_3892_45 <= _T_2797;
      end else begin
        _T_3892_45 <= _T_2594;
      end
    end
    if (_T_4005) begin
      if (_T_2891) begin
        _T_3892_46 <= _T_2798;
      end else begin
        _T_3892_46 <= _T_2595;
      end
    end
    if (_T_4006) begin
      if (_T_2891) begin
        _T_3892_47 <= _T_2799;
      end else begin
        _T_3892_47 <= _T_2596;
      end
    end
    if (_T_4007) begin
      if (_T_2891) begin
        _T_3892_48 <= _T_2800;
      end else begin
        _T_3892_48 <= _T_2597;
      end
    end
    if (_T_4008) begin
      if (_T_2891) begin
        _T_3892_49 <= _T_2801;
      end else begin
        _T_3892_49 <= _T_2598;
      end
    end
    if (_T_4009) begin
      if (_T_2891) begin
        _T_3892_50 <= _T_2802;
      end else begin
        _T_3892_50 <= _T_2599;
      end
    end
    if (_T_4010) begin
      if (_T_2891) begin
        _T_3892_51 <= _T_2803;
      end else begin
        _T_3892_51 <= _T_2600;
      end
    end
    if (_T_4011) begin
      if (_T_2891) begin
        _T_3892_52 <= _T_2804;
      end else begin
        _T_3892_52 <= _T_2601;
      end
    end
    if (_T_4012) begin
      if (_T_2891) begin
        _T_3892_53 <= _T_2805;
      end else begin
        _T_3892_53 <= _T_2602;
      end
    end
    if (_T_4013) begin
      if (_T_2891) begin
        _T_3892_54 <= _T_2806;
      end else begin
        _T_3892_54 <= _T_2603;
      end
    end
    if (_T_4014) begin
      if (_T_2891) begin
        _T_3892_55 <= _T_2807;
      end else begin
        _T_3892_55 <= _T_2604;
      end
    end
    if (_T_4015) begin
      if (_T_2891) begin
        _T_3892_56 <= _T_2808;
      end else begin
        _T_3892_56 <= _T_2605;
      end
    end
    if (_T_4016) begin
      if (_T_2891) begin
        _T_3892_57 <= _T_2809;
      end else begin
        _T_3892_57 <= _T_2606;
      end
    end
    if (_T_4017) begin
      if (_T_2891) begin
        _T_3892_58 <= _T_2810;
      end else begin
        _T_3892_58 <= _T_2607;
      end
    end
    if (_T_4018) begin
      if (_T_2891) begin
        _T_3892_59 <= _T_2811;
      end else begin
        _T_3892_59 <= _T_2608;
      end
    end
    if (_T_4019) begin
      if (_T_2891) begin
        _T_3892_60 <= _T_2812;
      end else begin
        _T_3892_60 <= _T_2609;
      end
    end
    if (_T_4020) begin
      if (_T_2891) begin
        _T_3892_61 <= _T_2813;
      end else begin
        _T_3892_61 <= _T_2610;
      end
    end
    if (_T_4021) begin
      if (_T_2891) begin
        _T_3892_62 <= _T_2814;
      end else begin
        _T_3892_62 <= _T_2611;
      end
    end
    if (_T_4022) begin
      if (_T_2891) begin
        _T_3892_63 <= _T_2815;
      end else begin
        _T_3892_63 <= _T_2612;
      end
    end
    if (_T_623) begin
      _T_4025 <= 1'h0;
    end else begin
      _T_4025 <= _T_3422;
    end
    if (_T_623) begin
      _T_4292_0 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_0 <= 1'h0;
        end else begin
          _T_4292_0 <= _T_3692_0;
        end
      end
    end
    if (_T_623) begin
      _T_4292_1 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_1 <= 1'h0;
        end else begin
          _T_4292_1 <= _T_3692_1;
        end
      end
    end
    if (_T_623) begin
      _T_4292_2 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_2 <= 1'h0;
        end else begin
          _T_4292_2 <= _T_3692_2;
        end
      end
    end
    if (_T_623) begin
      _T_4292_3 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_3 <= 1'h0;
        end else begin
          _T_4292_3 <= _T_3692_3;
        end
      end
    end
    if (_T_623) begin
      _T_4292_4 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_4 <= 1'h0;
        end else begin
          _T_4292_4 <= _T_3692_4;
        end
      end
    end
    if (_T_623) begin
      _T_4292_5 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_5 <= 1'h0;
        end else begin
          _T_4292_5 <= _T_3692_5;
        end
      end
    end
    if (_T_623) begin
      _T_4292_6 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_6 <= 1'h0;
        end else begin
          _T_4292_6 <= _T_3692_6;
        end
      end
    end
    if (_T_623) begin
      _T_4292_7 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_7 <= 1'h0;
        end else begin
          _T_4292_7 <= _T_3692_7;
        end
      end
    end
    if (_T_623) begin
      _T_4292_8 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_8 <= 1'h0;
        end else begin
          _T_4292_8 <= _T_3692_8;
        end
      end
    end
    if (_T_623) begin
      _T_4292_9 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_9 <= 1'h0;
        end else begin
          _T_4292_9 <= _T_3692_9;
        end
      end
    end
    if (_T_623) begin
      _T_4292_10 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_10 <= 1'h0;
        end else begin
          _T_4292_10 <= _T_3692_10;
        end
      end
    end
    if (_T_623) begin
      _T_4292_11 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_11 <= 1'h0;
        end else begin
          _T_4292_11 <= _T_3692_11;
        end
      end
    end
    if (_T_623) begin
      _T_4292_12 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_12 <= 1'h0;
        end else begin
          _T_4292_12 <= _T_3692_12;
        end
      end
    end
    if (_T_623) begin
      _T_4292_13 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_13 <= 1'h0;
        end else begin
          _T_4292_13 <= _T_3692_13;
        end
      end
    end
    if (_T_623) begin
      _T_4292_14 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_14 <= 1'h0;
        end else begin
          _T_4292_14 <= _T_3692_14;
        end
      end
    end
    if (_T_623) begin
      _T_4292_15 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_15 <= 1'h0;
        end else begin
          _T_4292_15 <= _T_3692_15;
        end
      end
    end
    if (_T_623) begin
      _T_4292_16 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_16 <= 1'h0;
        end else begin
          _T_4292_16 <= _T_3692_16;
        end
      end
    end
    if (_T_623) begin
      _T_4292_17 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_17 <= 1'h0;
        end else begin
          _T_4292_17 <= _T_3692_17;
        end
      end
    end
    if (_T_623) begin
      _T_4292_18 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_18 <= 1'h0;
        end else begin
          _T_4292_18 <= _T_3692_18;
        end
      end
    end
    if (_T_623) begin
      _T_4292_19 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_19 <= 1'h0;
        end else begin
          _T_4292_19 <= _T_3692_19;
        end
      end
    end
    if (_T_623) begin
      _T_4292_20 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_20 <= 1'h0;
        end else begin
          _T_4292_20 <= _T_3692_20;
        end
      end
    end
    if (_T_623) begin
      _T_4292_21 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_21 <= 1'h0;
        end else begin
          _T_4292_21 <= _T_3692_21;
        end
      end
    end
    if (_T_623) begin
      _T_4292_22 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_22 <= 1'h0;
        end else begin
          _T_4292_22 <= _T_3692_22;
        end
      end
    end
    if (_T_623) begin
      _T_4292_23 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_23 <= 1'h0;
        end else begin
          _T_4292_23 <= _T_3692_23;
        end
      end
    end
    if (_T_623) begin
      _T_4292_24 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_24 <= 1'h0;
        end else begin
          _T_4292_24 <= _T_3692_24;
        end
      end
    end
    if (_T_623) begin
      _T_4292_25 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_25 <= 1'h0;
        end else begin
          _T_4292_25 <= _T_3692_25;
        end
      end
    end
    if (_T_623) begin
      _T_4292_26 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_26 <= 1'h0;
        end else begin
          _T_4292_26 <= _T_3692_26;
        end
      end
    end
    if (_T_623) begin
      _T_4292_27 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_27 <= 1'h0;
        end else begin
          _T_4292_27 <= _T_3692_27;
        end
      end
    end
    if (_T_623) begin
      _T_4292_28 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_28 <= 1'h0;
        end else begin
          _T_4292_28 <= _T_3692_28;
        end
      end
    end
    if (_T_623) begin
      _T_4292_29 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_29 <= 1'h0;
        end else begin
          _T_4292_29 <= _T_3692_29;
        end
      end
    end
    if (_T_623) begin
      _T_4292_30 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_30 <= 1'h0;
        end else begin
          _T_4292_30 <= _T_3692_30;
        end
      end
    end
    if (_T_623) begin
      _T_4292_31 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_31 <= 1'h0;
        end else begin
          _T_4292_31 <= _T_3692_31;
        end
      end
    end
    if (_T_623) begin
      _T_4292_32 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_32 <= 1'h0;
        end else begin
          _T_4292_32 <= _T_3692_32;
        end
      end
    end
    if (_T_623) begin
      _T_4292_33 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_33 <= 1'h0;
        end else begin
          _T_4292_33 <= _T_3692_33;
        end
      end
    end
    if (_T_623) begin
      _T_4292_34 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_34 <= 1'h0;
        end else begin
          _T_4292_34 <= _T_3692_34;
        end
      end
    end
    if (_T_623) begin
      _T_4292_35 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_35 <= 1'h0;
        end else begin
          _T_4292_35 <= _T_3692_35;
        end
      end
    end
    if (_T_623) begin
      _T_4292_36 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_36 <= 1'h0;
        end else begin
          _T_4292_36 <= _T_3692_36;
        end
      end
    end
    if (_T_623) begin
      _T_4292_37 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_37 <= 1'h0;
        end else begin
          _T_4292_37 <= _T_3692_37;
        end
      end
    end
    if (_T_623) begin
      _T_4292_38 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_38 <= 1'h0;
        end else begin
          _T_4292_38 <= _T_3692_38;
        end
      end
    end
    if (_T_623) begin
      _T_4292_39 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_39 <= 1'h0;
        end else begin
          _T_4292_39 <= _T_3692_39;
        end
      end
    end
    if (_T_623) begin
      _T_4292_40 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_40 <= 1'h0;
        end else begin
          _T_4292_40 <= _T_3692_40;
        end
      end
    end
    if (_T_623) begin
      _T_4292_41 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_41 <= 1'h0;
        end else begin
          _T_4292_41 <= _T_3692_41;
        end
      end
    end
    if (_T_623) begin
      _T_4292_42 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_42 <= 1'h0;
        end else begin
          _T_4292_42 <= _T_3692_42;
        end
      end
    end
    if (_T_623) begin
      _T_4292_43 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_43 <= 1'h0;
        end else begin
          _T_4292_43 <= _T_3692_43;
        end
      end
    end
    if (_T_623) begin
      _T_4292_44 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_44 <= 1'h0;
        end else begin
          _T_4292_44 <= _T_3692_44;
        end
      end
    end
    if (_T_623) begin
      _T_4292_45 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_45 <= 1'h0;
        end else begin
          _T_4292_45 <= _T_3692_45;
        end
      end
    end
    if (_T_623) begin
      _T_4292_46 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_46 <= 1'h0;
        end else begin
          _T_4292_46 <= _T_3692_46;
        end
      end
    end
    if (_T_623) begin
      _T_4292_47 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_47 <= 1'h0;
        end else begin
          _T_4292_47 <= _T_3692_47;
        end
      end
    end
    if (_T_623) begin
      _T_4292_48 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_48 <= 1'h0;
        end else begin
          _T_4292_48 <= _T_3692_48;
        end
      end
    end
    if (_T_623) begin
      _T_4292_49 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_49 <= 1'h0;
        end else begin
          _T_4292_49 <= _T_3692_49;
        end
      end
    end
    if (_T_623) begin
      _T_4292_50 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_50 <= 1'h0;
        end else begin
          _T_4292_50 <= _T_3692_50;
        end
      end
    end
    if (_T_623) begin
      _T_4292_51 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_51 <= 1'h0;
        end else begin
          _T_4292_51 <= _T_3692_51;
        end
      end
    end
    if (_T_623) begin
      _T_4292_52 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_52 <= 1'h0;
        end else begin
          _T_4292_52 <= _T_3692_52;
        end
      end
    end
    if (_T_623) begin
      _T_4292_53 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_53 <= 1'h0;
        end else begin
          _T_4292_53 <= _T_3692_53;
        end
      end
    end
    if (_T_623) begin
      _T_4292_54 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_54 <= 1'h0;
        end else begin
          _T_4292_54 <= _T_3692_54;
        end
      end
    end
    if (_T_623) begin
      _T_4292_55 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_55 <= 1'h0;
        end else begin
          _T_4292_55 <= _T_3692_55;
        end
      end
    end
    if (_T_623) begin
      _T_4292_56 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_56 <= 1'h0;
        end else begin
          _T_4292_56 <= _T_3692_56;
        end
      end
    end
    if (_T_623) begin
      _T_4292_57 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_57 <= 1'h0;
        end else begin
          _T_4292_57 <= _T_3692_57;
        end
      end
    end
    if (_T_623) begin
      _T_4292_58 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_58 <= 1'h0;
        end else begin
          _T_4292_58 <= _T_3692_58;
        end
      end
    end
    if (_T_623) begin
      _T_4292_59 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_59 <= 1'h0;
        end else begin
          _T_4292_59 <= _T_3692_59;
        end
      end
    end
    if (_T_623) begin
      _T_4292_60 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_60 <= 1'h0;
        end else begin
          _T_4292_60 <= _T_3692_60;
        end
      end
    end
    if (_T_623) begin
      _T_4292_61 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_61 <= 1'h0;
        end else begin
          _T_4292_61 <= _T_3692_61;
        end
      end
    end
    if (_T_623) begin
      _T_4292_62 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_62 <= 1'h0;
        end else begin
          _T_4292_62 <= _T_3692_62;
        end
      end
    end
    if (_T_623) begin
      _T_4292_63 <= 1'h0;
    end else begin
      if (_T_4829) begin
        if (_T_4562) begin
          _T_4292_63 <= 1'h0;
        end else begin
          _T_4292_63 <= _T_3692_63;
        end
      end
    end
    if (_T_623) begin
      _T_4491 <= 9'h0;
    end else begin
      if (_T_3422) begin
        _T_4491 <= {{8'd0}, _T_3422};
      end
    end
    if (_T_4697_0) begin
      _T_4495_0 <= _T_3892_0;
    end
    if (_T_4697_1) begin
      _T_4495_1 <= _T_3892_1;
    end
    if (_T_4697_2) begin
      _T_4495_2 <= _T_3892_2;
    end
    if (_T_4697_3) begin
      _T_4495_3 <= _T_3892_3;
    end
    if (_T_4697_4) begin
      _T_4495_4 <= _T_3892_4;
    end
    if (_T_4697_5) begin
      _T_4495_5 <= _T_3892_5;
    end
    if (_T_4697_6) begin
      _T_4495_6 <= _T_3892_6;
    end
    if (_T_4697_7) begin
      _T_4495_7 <= _T_3892_7;
    end
    if (_T_4697_8) begin
      _T_4495_8 <= _T_3892_8;
    end
    if (_T_4697_9) begin
      _T_4495_9 <= _T_3892_9;
    end
    if (_T_4697_10) begin
      _T_4495_10 <= _T_3892_10;
    end
    if (_T_4697_11) begin
      _T_4495_11 <= _T_3892_11;
    end
    if (_T_4697_12) begin
      _T_4495_12 <= _T_3892_12;
    end
    if (_T_4697_13) begin
      _T_4495_13 <= _T_3892_13;
    end
    if (_T_4697_14) begin
      _T_4495_14 <= _T_3892_14;
    end
    if (_T_4697_15) begin
      _T_4495_15 <= _T_3892_15;
    end
    if (_T_4697_16) begin
      _T_4495_16 <= _T_3892_16;
    end
    if (_T_4697_17) begin
      _T_4495_17 <= _T_3892_17;
    end
    if (_T_4697_18) begin
      _T_4495_18 <= _T_3892_18;
    end
    if (_T_4697_19) begin
      _T_4495_19 <= _T_3892_19;
    end
    if (_T_4697_20) begin
      _T_4495_20 <= _T_3892_20;
    end
    if (_T_4697_21) begin
      _T_4495_21 <= _T_3892_21;
    end
    if (_T_4697_22) begin
      _T_4495_22 <= _T_3892_22;
    end
    if (_T_4697_23) begin
      _T_4495_23 <= _T_3892_23;
    end
    if (_T_4697_24) begin
      _T_4495_24 <= _T_3892_24;
    end
    if (_T_4697_25) begin
      _T_4495_25 <= _T_3892_25;
    end
    if (_T_4697_26) begin
      _T_4495_26 <= _T_3892_26;
    end
    if (_T_4697_27) begin
      _T_4495_27 <= _T_3892_27;
    end
    if (_T_4697_28) begin
      _T_4495_28 <= _T_3892_28;
    end
    if (_T_4697_29) begin
      _T_4495_29 <= _T_3892_29;
    end
    if (_T_4697_30) begin
      _T_4495_30 <= _T_3892_30;
    end
    if (_T_4697_31) begin
      _T_4495_31 <= _T_3892_31;
    end
    if (_T_4697_32) begin
      _T_4495_32 <= _T_3892_32;
    end
    if (_T_4697_33) begin
      _T_4495_33 <= _T_3892_33;
    end
    if (_T_4697_34) begin
      _T_4495_34 <= _T_3892_34;
    end
    if (_T_4697_35) begin
      _T_4495_35 <= _T_3892_35;
    end
    if (_T_4697_36) begin
      _T_4495_36 <= _T_3892_36;
    end
    if (_T_4697_37) begin
      _T_4495_37 <= _T_3892_37;
    end
    if (_T_4697_38) begin
      _T_4495_38 <= _T_3892_38;
    end
    if (_T_4697_39) begin
      _T_4495_39 <= _T_3892_39;
    end
    if (_T_4697_40) begin
      _T_4495_40 <= _T_3892_40;
    end
    if (_T_4697_41) begin
      _T_4495_41 <= _T_3892_41;
    end
    if (_T_4697_42) begin
      _T_4495_42 <= _T_3892_42;
    end
    if (_T_4697_43) begin
      _T_4495_43 <= _T_3892_43;
    end
    if (_T_4697_44) begin
      _T_4495_44 <= _T_3892_44;
    end
    if (_T_4697_45) begin
      _T_4495_45 <= _T_3892_45;
    end
    if (_T_4697_46) begin
      _T_4495_46 <= _T_3892_46;
    end
    if (_T_4697_47) begin
      _T_4495_47 <= _T_3892_47;
    end
    if (_T_4697_48) begin
      _T_4495_48 <= _T_3892_48;
    end
    if (_T_4697_49) begin
      _T_4495_49 <= _T_3892_49;
    end
    if (_T_4697_50) begin
      _T_4495_50 <= _T_3892_50;
    end
    if (_T_4697_51) begin
      _T_4495_51 <= _T_3892_51;
    end
    if (_T_4697_52) begin
      _T_4495_52 <= _T_3892_52;
    end
    if (_T_4697_53) begin
      _T_4495_53 <= _T_3892_53;
    end
    if (_T_4697_54) begin
      _T_4495_54 <= _T_3892_54;
    end
    if (_T_4697_55) begin
      _T_4495_55 <= _T_3892_55;
    end
    if (_T_4697_56) begin
      _T_4495_56 <= _T_3892_56;
    end
    if (_T_4697_57) begin
      _T_4495_57 <= _T_3892_57;
    end
    if (_T_4697_58) begin
      _T_4495_58 <= _T_3892_58;
    end
    if (_T_4697_59) begin
      _T_4495_59 <= _T_3892_59;
    end
    if (_T_4697_60) begin
      _T_4495_60 <= _T_3892_60;
    end
    if (_T_4697_61) begin
      _T_4495_61 <= _T_3892_61;
    end
    if (_T_4697_62) begin
      _T_4495_62 <= _T_3892_62;
    end
    if (_T_4697_63) begin
      _T_4495_63 <= _T_3892_63;
    end
    if (_T_623) begin
      _T_4832 <= 1'h0;
    end else begin
      _T_4832 <= _T_4025;
    end
    if (_T_623) begin
      _T_4838 <= 1'h0;
    end else begin
      _T_4838 <= _T_4025;
    end
    if (_T_623) begin
      _T_4841 <= 1'h0;
    end else begin
      _T_4841 <= _T_4025;
    end
    if (_T_623) begin
      _T_4845 <= 9'h0;
    end else begin
      if (_T_4843) begin
        if (_T_4833) begin
          _T_4845 <= 9'h0;
        end else begin
          _T_4845 <= _T_4491;
        end
      end
    end
    if (_T_623) begin
      _T_4849 <= 9'h0;
    end else begin
      if (_T_4843) begin
        if (_T_4833) begin
          _T_4849 <= 9'h0;
        end else begin
          _T_4849 <= _T_4491;
        end
      end
    end
    if (_T_623) begin
      _T_5117_0 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_0 <= _T_4292_0;
      end
    end
    if (_T_623) begin
      _T_5117_1 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_1 <= _T_4292_1;
      end
    end
    if (_T_623) begin
      _T_5117_2 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_2 <= _T_4292_2;
      end
    end
    if (_T_623) begin
      _T_5117_3 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_3 <= _T_4292_3;
      end
    end
    if (_T_623) begin
      _T_5117_4 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_4 <= _T_4292_4;
      end
    end
    if (_T_623) begin
      _T_5117_5 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_5 <= _T_4292_5;
      end
    end
    if (_T_623) begin
      _T_5117_6 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_6 <= _T_4292_6;
      end
    end
    if (_T_623) begin
      _T_5117_7 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_7 <= _T_4292_7;
      end
    end
    if (_T_623) begin
      _T_5117_8 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_8 <= _T_4292_8;
      end
    end
    if (_T_623) begin
      _T_5117_9 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_9 <= _T_4292_9;
      end
    end
    if (_T_623) begin
      _T_5117_10 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_10 <= _T_4292_10;
      end
    end
    if (_T_623) begin
      _T_5117_11 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_11 <= _T_4292_11;
      end
    end
    if (_T_623) begin
      _T_5117_12 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_12 <= _T_4292_12;
      end
    end
    if (_T_623) begin
      _T_5117_13 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_13 <= _T_4292_13;
      end
    end
    if (_T_623) begin
      _T_5117_14 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_14 <= _T_4292_14;
      end
    end
    if (_T_623) begin
      _T_5117_15 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_15 <= _T_4292_15;
      end
    end
    if (_T_623) begin
      _T_5117_16 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_16 <= _T_4292_16;
      end
    end
    if (_T_623) begin
      _T_5117_17 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_17 <= _T_4292_17;
      end
    end
    if (_T_623) begin
      _T_5117_18 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_18 <= _T_4292_18;
      end
    end
    if (_T_623) begin
      _T_5117_19 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_19 <= _T_4292_19;
      end
    end
    if (_T_623) begin
      _T_5117_20 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_20 <= _T_4292_20;
      end
    end
    if (_T_623) begin
      _T_5117_21 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_21 <= _T_4292_21;
      end
    end
    if (_T_623) begin
      _T_5117_22 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_22 <= _T_4292_22;
      end
    end
    if (_T_623) begin
      _T_5117_23 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_23 <= _T_4292_23;
      end
    end
    if (_T_623) begin
      _T_5117_24 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_24 <= _T_4292_24;
      end
    end
    if (_T_623) begin
      _T_5117_25 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_25 <= _T_4292_25;
      end
    end
    if (_T_623) begin
      _T_5117_26 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_26 <= _T_4292_26;
      end
    end
    if (_T_623) begin
      _T_5117_27 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_27 <= _T_4292_27;
      end
    end
    if (_T_623) begin
      _T_5117_28 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_28 <= _T_4292_28;
      end
    end
    if (_T_623) begin
      _T_5117_29 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_29 <= _T_4292_29;
      end
    end
    if (_T_623) begin
      _T_5117_30 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_30 <= _T_4292_30;
      end
    end
    if (_T_623) begin
      _T_5117_31 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_31 <= _T_4292_31;
      end
    end
    if (_T_623) begin
      _T_5117_32 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_32 <= _T_4292_32;
      end
    end
    if (_T_623) begin
      _T_5117_33 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_33 <= _T_4292_33;
      end
    end
    if (_T_623) begin
      _T_5117_34 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_34 <= _T_4292_34;
      end
    end
    if (_T_623) begin
      _T_5117_35 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_35 <= _T_4292_35;
      end
    end
    if (_T_623) begin
      _T_5117_36 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_36 <= _T_4292_36;
      end
    end
    if (_T_623) begin
      _T_5117_37 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_37 <= _T_4292_37;
      end
    end
    if (_T_623) begin
      _T_5117_38 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_38 <= _T_4292_38;
      end
    end
    if (_T_623) begin
      _T_5117_39 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_39 <= _T_4292_39;
      end
    end
    if (_T_623) begin
      _T_5117_40 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_40 <= _T_4292_40;
      end
    end
    if (_T_623) begin
      _T_5117_41 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_41 <= _T_4292_41;
      end
    end
    if (_T_623) begin
      _T_5117_42 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_42 <= _T_4292_42;
      end
    end
    if (_T_623) begin
      _T_5117_43 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_43 <= _T_4292_43;
      end
    end
    if (_T_623) begin
      _T_5117_44 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_44 <= _T_4292_44;
      end
    end
    if (_T_623) begin
      _T_5117_45 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_45 <= _T_4292_45;
      end
    end
    if (_T_623) begin
      _T_5117_46 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_46 <= _T_4292_46;
      end
    end
    if (_T_623) begin
      _T_5117_47 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_47 <= _T_4292_47;
      end
    end
    if (_T_623) begin
      _T_5117_48 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_48 <= _T_4292_48;
      end
    end
    if (_T_623) begin
      _T_5117_49 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_49 <= _T_4292_49;
      end
    end
    if (_T_623) begin
      _T_5117_50 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_50 <= _T_4292_50;
      end
    end
    if (_T_623) begin
      _T_5117_51 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_51 <= _T_4292_51;
      end
    end
    if (_T_623) begin
      _T_5117_52 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_52 <= _T_4292_52;
      end
    end
    if (_T_623) begin
      _T_5117_53 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_53 <= _T_4292_53;
      end
    end
    if (_T_623) begin
      _T_5117_54 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_54 <= _T_4292_54;
      end
    end
    if (_T_623) begin
      _T_5117_55 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_55 <= _T_4292_55;
      end
    end
    if (_T_623) begin
      _T_5117_56 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_56 <= _T_4292_56;
      end
    end
    if (_T_623) begin
      _T_5117_57 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_57 <= _T_4292_57;
      end
    end
    if (_T_623) begin
      _T_5117_58 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_58 <= _T_4292_58;
      end
    end
    if (_T_623) begin
      _T_5117_59 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_59 <= _T_4292_59;
      end
    end
    if (_T_623) begin
      _T_5117_60 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_60 <= _T_4292_60;
      end
    end
    if (_T_623) begin
      _T_5117_61 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_61 <= _T_4292_61;
      end
    end
    if (_T_623) begin
      _T_5117_62 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_62 <= _T_4292_62;
      end
    end
    if (_T_623) begin
      _T_5117_63 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5117_63 <= _T_4292_63;
      end
    end
    if (_T_623) begin
      _T_5581_0 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_0 <= _T_4292_0;
      end
    end
    if (_T_623) begin
      _T_5581_1 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_1 <= _T_4292_1;
      end
    end
    if (_T_623) begin
      _T_5581_2 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_2 <= _T_4292_2;
      end
    end
    if (_T_623) begin
      _T_5581_3 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_3 <= _T_4292_3;
      end
    end
    if (_T_623) begin
      _T_5581_4 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_4 <= _T_4292_4;
      end
    end
    if (_T_623) begin
      _T_5581_5 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_5 <= _T_4292_5;
      end
    end
    if (_T_623) begin
      _T_5581_6 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_6 <= _T_4292_6;
      end
    end
    if (_T_623) begin
      _T_5581_7 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_7 <= _T_4292_7;
      end
    end
    if (_T_623) begin
      _T_5581_8 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_8 <= _T_4292_8;
      end
    end
    if (_T_623) begin
      _T_5581_9 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_9 <= _T_4292_9;
      end
    end
    if (_T_623) begin
      _T_5581_10 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_10 <= _T_4292_10;
      end
    end
    if (_T_623) begin
      _T_5581_11 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_11 <= _T_4292_11;
      end
    end
    if (_T_623) begin
      _T_5581_12 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_12 <= _T_4292_12;
      end
    end
    if (_T_623) begin
      _T_5581_13 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_13 <= _T_4292_13;
      end
    end
    if (_T_623) begin
      _T_5581_14 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_14 <= _T_4292_14;
      end
    end
    if (_T_623) begin
      _T_5581_15 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_15 <= _T_4292_15;
      end
    end
    if (_T_623) begin
      _T_5581_16 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_16 <= _T_4292_16;
      end
    end
    if (_T_623) begin
      _T_5581_17 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_17 <= _T_4292_17;
      end
    end
    if (_T_623) begin
      _T_5581_18 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_18 <= _T_4292_18;
      end
    end
    if (_T_623) begin
      _T_5581_19 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_19 <= _T_4292_19;
      end
    end
    if (_T_623) begin
      _T_5581_20 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_20 <= _T_4292_20;
      end
    end
    if (_T_623) begin
      _T_5581_21 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_21 <= _T_4292_21;
      end
    end
    if (_T_623) begin
      _T_5581_22 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_22 <= _T_4292_22;
      end
    end
    if (_T_623) begin
      _T_5581_23 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_23 <= _T_4292_23;
      end
    end
    if (_T_623) begin
      _T_5581_24 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_24 <= _T_4292_24;
      end
    end
    if (_T_623) begin
      _T_5581_25 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_25 <= _T_4292_25;
      end
    end
    if (_T_623) begin
      _T_5581_26 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_26 <= _T_4292_26;
      end
    end
    if (_T_623) begin
      _T_5581_27 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_27 <= _T_4292_27;
      end
    end
    if (_T_623) begin
      _T_5581_28 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_28 <= _T_4292_28;
      end
    end
    if (_T_623) begin
      _T_5581_29 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_29 <= _T_4292_29;
      end
    end
    if (_T_623) begin
      _T_5581_30 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_30 <= _T_4292_30;
      end
    end
    if (_T_623) begin
      _T_5581_31 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_31 <= _T_4292_31;
      end
    end
    if (_T_623) begin
      _T_5581_32 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_32 <= _T_4292_32;
      end
    end
    if (_T_623) begin
      _T_5581_33 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_33 <= _T_4292_33;
      end
    end
    if (_T_623) begin
      _T_5581_34 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_34 <= _T_4292_34;
      end
    end
    if (_T_623) begin
      _T_5581_35 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_35 <= _T_4292_35;
      end
    end
    if (_T_623) begin
      _T_5581_36 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_36 <= _T_4292_36;
      end
    end
    if (_T_623) begin
      _T_5581_37 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_37 <= _T_4292_37;
      end
    end
    if (_T_623) begin
      _T_5581_38 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_38 <= _T_4292_38;
      end
    end
    if (_T_623) begin
      _T_5581_39 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_39 <= _T_4292_39;
      end
    end
    if (_T_623) begin
      _T_5581_40 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_40 <= _T_4292_40;
      end
    end
    if (_T_623) begin
      _T_5581_41 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_41 <= _T_4292_41;
      end
    end
    if (_T_623) begin
      _T_5581_42 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_42 <= _T_4292_42;
      end
    end
    if (_T_623) begin
      _T_5581_43 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_43 <= _T_4292_43;
      end
    end
    if (_T_623) begin
      _T_5581_44 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_44 <= _T_4292_44;
      end
    end
    if (_T_623) begin
      _T_5581_45 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_45 <= _T_4292_45;
      end
    end
    if (_T_623) begin
      _T_5581_46 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_46 <= _T_4292_46;
      end
    end
    if (_T_623) begin
      _T_5581_47 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_47 <= _T_4292_47;
      end
    end
    if (_T_623) begin
      _T_5581_48 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_48 <= _T_4292_48;
      end
    end
    if (_T_623) begin
      _T_5581_49 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_49 <= _T_4292_49;
      end
    end
    if (_T_623) begin
      _T_5581_50 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_50 <= _T_4292_50;
      end
    end
    if (_T_623) begin
      _T_5581_51 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_51 <= _T_4292_51;
      end
    end
    if (_T_623) begin
      _T_5581_52 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_52 <= _T_4292_52;
      end
    end
    if (_T_623) begin
      _T_5581_53 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_53 <= _T_4292_53;
      end
    end
    if (_T_623) begin
      _T_5581_54 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_54 <= _T_4292_54;
      end
    end
    if (_T_623) begin
      _T_5581_55 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_55 <= _T_4292_55;
      end
    end
    if (_T_623) begin
      _T_5581_56 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_56 <= _T_4292_56;
      end
    end
    if (_T_623) begin
      _T_5581_57 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_57 <= _T_4292_57;
      end
    end
    if (_T_623) begin
      _T_5581_58 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_58 <= _T_4292_58;
      end
    end
    if (_T_623) begin
      _T_5581_59 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_59 <= _T_4292_59;
      end
    end
    if (_T_623) begin
      _T_5581_60 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_60 <= _T_4292_60;
      end
    end
    if (_T_623) begin
      _T_5581_61 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_61 <= _T_4292_61;
      end
    end
    if (_T_623) begin
      _T_5581_62 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_62 <= _T_4292_62;
      end
    end
    if (_T_623) begin
      _T_5581_63 <= 1'h0;
    end else begin
      if (_T_4843) begin
        _T_5581_63 <= _T_4292_63;
      end
    end
    if (_T_4292_0) begin
      _T_5779 <= _T_4495_0;
    end
    if (_T_4292_0) begin
      _T_5781 <= _T_4495_0;
    end
    if (_T_4292_1) begin
      _T_5783 <= _T_4495_1;
    end
    if (_T_4292_1) begin
      _T_5785 <= _T_4495_1;
    end
    if (_T_4292_2) begin
      _T_5787 <= _T_4495_2;
    end
    if (_T_4292_2) begin
      _T_5789 <= _T_4495_2;
    end
    if (_T_4292_3) begin
      _T_5791 <= _T_4495_3;
    end
    if (_T_4292_3) begin
      _T_5793 <= _T_4495_3;
    end
    if (_T_4292_4) begin
      _T_5795 <= _T_4495_4;
    end
    if (_T_4292_4) begin
      _T_5797 <= _T_4495_4;
    end
    if (_T_4292_5) begin
      _T_5799 <= _T_4495_5;
    end
    if (_T_4292_5) begin
      _T_5801 <= _T_4495_5;
    end
    if (_T_4292_6) begin
      _T_5803 <= _T_4495_6;
    end
    if (_T_4292_6) begin
      _T_5805 <= _T_4495_6;
    end
    if (_T_4292_7) begin
      _T_5807 <= _T_4495_7;
    end
    if (_T_4292_7) begin
      _T_5809 <= _T_4495_7;
    end
    if (_T_4292_8) begin
      _T_5811 <= _T_4495_8;
    end
    if (_T_4292_8) begin
      _T_5813 <= _T_4495_8;
    end
    if (_T_4292_9) begin
      _T_5815 <= _T_4495_9;
    end
    if (_T_4292_9) begin
      _T_5817 <= _T_4495_9;
    end
    if (_T_4292_10) begin
      _T_5819 <= _T_4495_10;
    end
    if (_T_4292_10) begin
      _T_5821 <= _T_4495_10;
    end
    if (_T_4292_11) begin
      _T_5823 <= _T_4495_11;
    end
    if (_T_4292_11) begin
      _T_5825 <= _T_4495_11;
    end
    if (_T_4292_12) begin
      _T_5827 <= _T_4495_12;
    end
    if (_T_4292_12) begin
      _T_5829 <= _T_4495_12;
    end
    if (_T_4292_13) begin
      _T_5831 <= _T_4495_13;
    end
    if (_T_4292_13) begin
      _T_5833 <= _T_4495_13;
    end
    if (_T_4292_14) begin
      _T_5835 <= _T_4495_14;
    end
    if (_T_4292_14) begin
      _T_5837 <= _T_4495_14;
    end
    if (_T_4292_15) begin
      _T_5839 <= _T_4495_15;
    end
    if (_T_4292_15) begin
      _T_5841 <= _T_4495_15;
    end
    if (_T_4292_16) begin
      _T_5843 <= _T_4495_16;
    end
    if (_T_4292_16) begin
      _T_5845 <= _T_4495_16;
    end
    if (_T_4292_17) begin
      _T_5847 <= _T_4495_17;
    end
    if (_T_4292_17) begin
      _T_5849 <= _T_4495_17;
    end
    if (_T_4292_18) begin
      _T_5851 <= _T_4495_18;
    end
    if (_T_4292_18) begin
      _T_5853 <= _T_4495_18;
    end
    if (_T_4292_19) begin
      _T_5855 <= _T_4495_19;
    end
    if (_T_4292_19) begin
      _T_5857 <= _T_4495_19;
    end
    if (_T_4292_20) begin
      _T_5859 <= _T_4495_20;
    end
    if (_T_4292_20) begin
      _T_5861 <= _T_4495_20;
    end
    if (_T_4292_21) begin
      _T_5863 <= _T_4495_21;
    end
    if (_T_4292_21) begin
      _T_5865 <= _T_4495_21;
    end
    if (_T_4292_22) begin
      _T_5867 <= _T_4495_22;
    end
    if (_T_4292_22) begin
      _T_5869 <= _T_4495_22;
    end
    if (_T_4292_23) begin
      _T_5871 <= _T_4495_23;
    end
    if (_T_4292_23) begin
      _T_5873 <= _T_4495_23;
    end
    if (_T_4292_24) begin
      _T_5875 <= _T_4495_24;
    end
    if (_T_4292_24) begin
      _T_5877 <= _T_4495_24;
    end
    if (_T_4292_25) begin
      _T_5879 <= _T_4495_25;
    end
    if (_T_4292_25) begin
      _T_5881 <= _T_4495_25;
    end
    if (_T_4292_26) begin
      _T_5883 <= _T_4495_26;
    end
    if (_T_4292_26) begin
      _T_5885 <= _T_4495_26;
    end
    if (_T_4292_27) begin
      _T_5887 <= _T_4495_27;
    end
    if (_T_4292_27) begin
      _T_5889 <= _T_4495_27;
    end
    if (_T_4292_28) begin
      _T_5891 <= _T_4495_28;
    end
    if (_T_4292_28) begin
      _T_5893 <= _T_4495_28;
    end
    if (_T_4292_29) begin
      _T_5895 <= _T_4495_29;
    end
    if (_T_4292_29) begin
      _T_5897 <= _T_4495_29;
    end
    if (_T_4292_30) begin
      _T_5899 <= _T_4495_30;
    end
    if (_T_4292_30) begin
      _T_5901 <= _T_4495_30;
    end
    if (_T_4292_31) begin
      _T_5903 <= _T_4495_31;
    end
    if (_T_4292_31) begin
      _T_5905 <= _T_4495_31;
    end
    if (_T_4292_32) begin
      _T_5907 <= _T_4495_32;
    end
    if (_T_4292_32) begin
      _T_5909 <= _T_4495_32;
    end
    if (_T_4292_33) begin
      _T_5911 <= _T_4495_33;
    end
    if (_T_4292_33) begin
      _T_5913 <= _T_4495_33;
    end
    if (_T_4292_34) begin
      _T_5915 <= _T_4495_34;
    end
    if (_T_4292_34) begin
      _T_5917 <= _T_4495_34;
    end
    if (_T_4292_35) begin
      _T_5919 <= _T_4495_35;
    end
    if (_T_4292_35) begin
      _T_5921 <= _T_4495_35;
    end
    if (_T_4292_36) begin
      _T_5923 <= _T_4495_36;
    end
    if (_T_4292_36) begin
      _T_5925 <= _T_4495_36;
    end
    if (_T_4292_37) begin
      _T_5927 <= _T_4495_37;
    end
    if (_T_4292_37) begin
      _T_5929 <= _T_4495_37;
    end
    if (_T_4292_38) begin
      _T_5931 <= _T_4495_38;
    end
    if (_T_4292_38) begin
      _T_5933 <= _T_4495_38;
    end
    if (_T_4292_39) begin
      _T_5935 <= _T_4495_39;
    end
    if (_T_4292_39) begin
      _T_5937 <= _T_4495_39;
    end
    if (_T_4292_40) begin
      _T_5939 <= _T_4495_40;
    end
    if (_T_4292_40) begin
      _T_5941 <= _T_4495_40;
    end
    if (_T_4292_41) begin
      _T_5943 <= _T_4495_41;
    end
    if (_T_4292_41) begin
      _T_5945 <= _T_4495_41;
    end
    if (_T_4292_42) begin
      _T_5947 <= _T_4495_42;
    end
    if (_T_4292_42) begin
      _T_5949 <= _T_4495_42;
    end
    if (_T_4292_43) begin
      _T_5951 <= _T_4495_43;
    end
    if (_T_4292_43) begin
      _T_5953 <= _T_4495_43;
    end
    if (_T_4292_44) begin
      _T_5955 <= _T_4495_44;
    end
    if (_T_4292_44) begin
      _T_5957 <= _T_4495_44;
    end
    if (_T_4292_45) begin
      _T_5959 <= _T_4495_45;
    end
    if (_T_4292_45) begin
      _T_5961 <= _T_4495_45;
    end
    if (_T_4292_46) begin
      _T_5963 <= _T_4495_46;
    end
    if (_T_4292_46) begin
      _T_5965 <= _T_4495_46;
    end
    if (_T_4292_47) begin
      _T_5967 <= _T_4495_47;
    end
    if (_T_4292_47) begin
      _T_5969 <= _T_4495_47;
    end
    if (_T_4292_48) begin
      _T_5971 <= _T_4495_48;
    end
    if (_T_4292_48) begin
      _T_5973 <= _T_4495_48;
    end
    if (_T_4292_49) begin
      _T_5975 <= _T_4495_49;
    end
    if (_T_4292_49) begin
      _T_5977 <= _T_4495_49;
    end
    if (_T_4292_50) begin
      _T_5979 <= _T_4495_50;
    end
    if (_T_4292_50) begin
      _T_5981 <= _T_4495_50;
    end
    if (_T_4292_51) begin
      _T_5983 <= _T_4495_51;
    end
    if (_T_4292_51) begin
      _T_5985 <= _T_4495_51;
    end
    if (_T_4292_52) begin
      _T_5987 <= _T_4495_52;
    end
    if (_T_4292_52) begin
      _T_5989 <= _T_4495_52;
    end
    if (_T_4292_53) begin
      _T_5991 <= _T_4495_53;
    end
    if (_T_4292_53) begin
      _T_5993 <= _T_4495_53;
    end
    if (_T_4292_54) begin
      _T_5995 <= _T_4495_54;
    end
    if (_T_4292_54) begin
      _T_5997 <= _T_4495_54;
    end
    if (_T_4292_55) begin
      _T_5999 <= _T_4495_55;
    end
    if (_T_4292_55) begin
      _T_6001 <= _T_4495_55;
    end
    if (_T_4292_56) begin
      _T_6003 <= _T_4495_56;
    end
    if (_T_4292_56) begin
      _T_6005 <= _T_4495_56;
    end
    if (_T_4292_57) begin
      _T_6007 <= _T_4495_57;
    end
    if (_T_4292_57) begin
      _T_6009 <= _T_4495_57;
    end
    if (_T_4292_58) begin
      _T_6011 <= _T_4495_58;
    end
    if (_T_4292_58) begin
      _T_6013 <= _T_4495_58;
    end
    if (_T_4292_59) begin
      _T_6015 <= _T_4495_59;
    end
    if (_T_4292_59) begin
      _T_6017 <= _T_4495_59;
    end
    if (_T_4292_60) begin
      _T_6019 <= _T_4495_60;
    end
    if (_T_4292_60) begin
      _T_6021 <= _T_4495_60;
    end
    if (_T_4292_61) begin
      _T_6023 <= _T_4495_61;
    end
    if (_T_4292_61) begin
      _T_6025 <= _T_4495_61;
    end
    if (_T_4292_62) begin
      _T_6027 <= _T_4495_62;
    end
    if (_T_4292_62) begin
      _T_6029 <= _T_4495_62;
    end
    if (_T_4292_63) begin
      _T_6031 <= _T_4495_63;
    end
    if (_T_4292_63) begin
      _T_6033 <= _T_4495_63;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (_T_623) begin
      _T_1079 <= 15'h0;
    end else begin
      if (_T_1151) begin
        if (io_sc2cdma_dat_pending_req) begin
          _T_1079 <= 15'h0;
        end else begin
          if (_T_1122) begin
            _T_1079 <= _T_1115;
          end else begin
            _T_1079 <= _T_1106;
          end
        end
      end
    end
  end
endmodule

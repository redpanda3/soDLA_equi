module NV_soDLA_CSC_dl_for_check( // @[:@3.2]
  input          nvdla_core_clk, // @[:@6.4]
  input          nvdla_core_ng_clk, // @[:@6.4]
  input          nvdla_core_rstn, // @[:@6.4]
  input  [1:0]   sc_state, // @[:@6.4]
  input          sg2dl_reuse_rls, // @[:@6.4]
  input          sg2dl_pvld, // @[:@6.4]
  input  [30:0]  sg2dl_pd, // @[:@6.4]
  input          cdma2sc_dat_updt, // @[:@6.4]
  input  [14:0]  cdma2sc_dat_entries, // @[:@6.4]
  input  [13:0]  cdma2sc_dat_slices, // @[:@6.4]
  input          sc2cdma_dat_pending_req, // @[:@6.4]
  output         sc2cdma_dat_updt, // @[:@6.4]
  output [14:0]  sc2cdma_dat_entries, // @[:@6.4]
  output [13:0]  sc2cdma_dat_slices, // @[:@6.4]
  output         sc2buf_dat_rd_en, // @[:@6.4]
  output [12:0]  sc2buf_dat_rd_addr, // @[:@6.4]
  input          sc2buf_dat_rd_valid, // @[:@6.4]
  input  [511:0] sc2buf_dat_rd_data, // @[:@6.4]
  output         sc2mac_dat_a_pvld, // @[:@6.4]
  output [63:0]  sc2mac_dat_a_mask, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data0, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data1, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data2, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data3, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data4, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data5, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data6, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data7, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data8, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data9, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data10, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data11, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data12, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data13, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data14, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data15, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data16, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data17, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data18, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data19, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data20, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data21, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data22, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data23, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data24, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data25, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data26, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data27, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data28, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data29, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data30, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data31, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data32, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data33, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data34, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data35, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data36, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data37, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data38, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data39, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data40, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data41, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data42, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data43, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data44, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data45, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data46, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data47, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data48, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data49, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data50, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data51, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data52, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data53, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data54, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data55, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data56, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data57, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data58, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data59, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data60, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data61, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data62, // @[:@6.4]
  output [7:0]   sc2mac_dat_a_data63, // @[:@6.4]
  output [8:0]   sc2mac_dat_a_pd, // @[:@6.4]
  output         sc2mac_dat_b_pvld, // @[:@6.4]
  output [63:0]  sc2mac_dat_b_mask, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data0, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data1, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data2, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data3, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data4, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data5, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data6, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data7, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data8, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data9, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data10, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data11, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data12, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data13, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data14, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data15, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data16, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data17, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data18, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data19, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data20, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data21, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data22, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data23, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data24, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data25, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data26, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data27, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data28, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data29, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data30, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data31, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data32, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data33, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data34, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data35, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data36, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data37, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data38, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data39, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data40, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data41, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data42, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data43, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data44, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data45, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data46, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data47, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data48, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data49, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data50, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data51, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data52, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data53, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data54, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data55, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data56, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data57, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data58, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data59, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data60, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data61, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data62, // @[:@6.4]
  output [7:0]   sc2mac_dat_b_data63, // @[:@6.4]
  output [8:0]   sc2mac_dat_b_pd, // @[:@6.4]
  input          reg2dp_op_en, // @[:@6.4]
  input          reg2dp_conv_mode, // @[:@6.4]
  input  [4:0]   reg2dp_batches, // @[:@6.4]
  input  [1:0]   reg2dp_proc_precision, // @[:@6.4]
  input          reg2dp_datain_format, // @[:@6.4]
  input          reg2dp_skip_data_rls, // @[:@6.4]
  input  [12:0]  reg2dp_datain_channel_ext, // @[:@6.4]
  input  [12:0]  reg2dp_datain_height_ext, // @[:@6.4]
  input  [12:0]  reg2dp_datain_width_ext, // @[:@6.4]
  input  [1:0]   reg2dp_y_extension, // @[:@6.4]
  input  [12:0]  reg2dp_weight_channel_ext, // @[:@6.4]
  input  [13:0]  reg2dp_entries, // @[:@6.4]
  input  [12:0]  reg2dp_dataout_width, // @[:@6.4]
  input  [11:0]  reg2dp_rls_slices, // @[:@6.4]
  input  [2:0]   reg2dp_conv_x_stride_ext, // @[:@6.4]
  input  [2:0]   reg2dp_conv_y_stride_ext, // @[:@6.4]
  input  [4:0]   reg2dp_x_dilation_ext, // @[:@6.4]
  input  [4:0]   reg2dp_y_dilation_ext, // @[:@6.4]
  input  [4:0]   reg2dp_pad_left, // @[:@6.4]
  input  [4:0]   reg2dp_pad_top, // @[:@6.4]
  input  [15:0]  reg2dp_pad_value, // @[:@6.4]
  input  [4:0]   reg2dp_data_bank, // @[:@6.4]
  input  [1:0]   reg2dp_pra_truncate, // @[:@6.4]
  output         slcg_wg_en // @[:@6.4]
);
  wire  _T_337; // @[NV_NVDLA_CSC_dl_for_check.scala 95:38:@8.4]
  wire  is_sg_idle; // @[NV_NVDLA_CSC_dl_for_check.scala 99:31:@9.4]
  wire  is_sg_done; // @[NV_NVDLA_CSC_dl_for_check.scala 101:31:@11.4]
  wire  layer_st; // @[NV_NVDLA_CSC_dl_for_check.scala 108:32:@14.4]
  wire  is_conv; // @[NV_NVDLA_CSC_dl_for_check.scala 110:35:@16.4]
  wire  is_img; // @[NV_NVDLA_CSC_dl_for_check.scala 111:22:@17.4]
  wire [6:0] _T_346; // @[NV_NVDLA_CSC_dl_for_check.scala 118:53:@18.4]
  wire [6:0] _T_348; // @[NV_NVDLA_CSC_dl_for_check.scala 118:24:@19.4]
  wire [2:0] sub_h_total_w; // @[NV_NVDLA_CSC_dl_for_check.scala 118:100:@20.4]
  wire [2:0] sub_h_cmp_w; // @[NV_NVDLA_CSC_dl_for_check.scala 119:22:@21.4]
  wire [3:0] _T_351; // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@22.4]
  wire [3:0] dataout_w_init; // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@23.4]
  wire [3:0] conv_x_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 121:51:@24.4]
  wire [1:0] _T_353; // @[NV_NVDLA_CSC_dl_for_check.scala 122:62:@25.4]
  wire [5:0] _T_356; // @[Cat.scala 30:58:@26.4]
  wire [4:0] _T_359; // @[Cat.scala 30:58:@27.4]
  wire [4:0] _GEN_671; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  wire [5:0] _T_360; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  wire  _T_361; // @[Mux.scala 46:19:@29.4]
  wire [5:0] _T_362; // @[Mux.scala 46:16:@30.4]
  wire  _T_363; // @[Mux.scala 46:19:@31.4]
  wire [5:0] pixel_x_stride_w; // @[Mux.scala 46:16:@32.4]
  wire  _T_365; // @[NV_NVDLA_CSC_dl_for_check.scala 126:88:@33.4]
  wire [5:0] _T_371; // @[NV_NVDLA_CSC_dl_for_check.scala 126:172:@35.4]
  wire [5:0] _T_372; // @[NV_NVDLA_CSC_dl_for_check.scala 126:58:@36.4]
  wire [6:0] _T_375; // @[Cat.scala 30:58:@37.4]
  wire [6:0] _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  wire [7:0] _T_376; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  wire [6:0] _T_377; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@39.4]
  wire [6:0] _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  wire [7:0] _T_379; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  wire [6:0] _T_380; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@42.4]
  wire [6:0] _T_383; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@44.4]
  wire [5:0] _T_384; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@45.4]
  wire  _T_385; // @[Mux.scala 46:19:@46.4]
  wire [5:0] _T_386; // @[Mux.scala 46:16:@47.4]
  wire  _T_387; // @[Mux.scala 46:19:@48.4]
  wire [6:0] pixel_x_init_w; // @[Mux.scala 46:16:@49.4]
  wire [6:0] pixel_x_init_offset_w; // @[NV_NVDLA_CSC_dl_for_check.scala 129:80:@51.4]
  wire [7:0] _T_392; // @[Cat.scala 30:58:@52.4]
  wire [6:0] _T_397; // @[Mux.scala 46:16:@55.4]
  wire [7:0] pixel_x_add_w; // @[Mux.scala 46:16:@57.4]
  wire [11:0] pixel_ch_stride_w; // @[Cat.scala 30:58:@58.4]
  wire [3:0] conv_y_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 139:52:@59.4]
  wire [5:0] _T_403; // @[NV_NVDLA_CSC_dl_for_check.scala 140:60:@60.4]
  wire [5:0] x_dilate_w; // @[NV_NVDLA_CSC_dl_for_check.scala 140:21:@61.4]
  wire [5:0] _T_406; // @[NV_NVDLA_CSC_dl_for_check.scala 141:60:@62.4]
  wire [5:0] y_dilate_w; // @[NV_NVDLA_CSC_dl_for_check.scala 141:21:@63.4]
  reg  layer_st_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 143:26:@64.4]
  reg [31:0] _RAND_0;
  reg [5:0] data_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 144:25:@66.4]
  reg [31:0] _RAND_1;
  reg [13:0] rls_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 145:25:@68.4]
  reg [31:0] _RAND_2;
  reg [13:0] h_offset_slice; // @[NV_NVDLA_CSC_dl_for_check.scala 146:29:@70.4]
  reg [31:0] _RAND_3;
  reg [14:0] entries; // @[NV_NVDLA_CSC_dl_for_check.scala 147:22:@72.4]
  reg [31:0] _RAND_4;
  reg [14:0] entries_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 148:28:@74.4]
  reg [31:0] _RAND_5;
  reg [12:0] dataout_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 149:32:@76.4]
  reg [31:0] _RAND_6;
  reg [14:0] rls_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 151:26:@80.4]
  reg [31:0] _RAND_7;
  reg [11:0] h_bias_0_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 152:30:@82.4]
  reg [31:0] _RAND_8;
  reg [11:0] h_bias_1_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 153:30:@84.4]
  reg [31:0] _RAND_9;
  reg [13:0] slice_left; // @[NV_NVDLA_CSC_dl_for_check.scala 154:25:@86.4]
  reg [31:0] _RAND_10;
  wire [14:0] entries_single_w; // @[NV_NVDLA_CSC_dl_for_check.scala 157:43:@87.4]
  wire [20:0] _T_477; // @[NV_NVDLA_CSC_dl_for_check.scala 158:41:@89.4]
  wire [14:0] entries_batch_w; // @[NV_NVDLA_CSC_dl_for_check.scala 158:56:@90.4]
  wire [11:0] h_offset_slice_w; // @[NV_NVDLA_CSC_dl_for_check.scala 160:37:@91.4]
  wire [14:0] _GEN_674; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  wire [20:0] _T_478; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  wire [11:0] h_bias_0_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 161:47:@93.4]
  wire [14:0] _GEN_675; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  wire [28:0] _T_479; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  wire [11:0] h_bias_1_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 162:51:@95.4]
  wire [12:0] rls_slices_w; // @[NV_NVDLA_CSC_dl_for_check.scala 163:41:@96.4]
  wire [13:0] _T_482; // @[NV_NVDLA_CSC_dl_for_check.scala 164:77:@97.4]
  wire [12:0] _GEN_676; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@98.4]
  wire [13:0] _T_483; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@98.4]
  wire [13:0] _T_484; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@99.4]
  wire [13:0] slice_left_w; // @[NV_NVDLA_CSC_dl_for_check.scala 164:23:@100.4]
  wire [13:0] slices_oprand; // @[NV_NVDLA_CSC_dl_for_check.scala 165:24:@101.4]
  wire [14:0] _GEN_677; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@102.4]
  wire [28:0] _T_485; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@102.4]
  wire [14:0] slice_entries_w; // @[NV_NVDLA_CSC_dl_for_check.scala 166:54:@103.4]
  reg [33:0] is_img_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 171:24:@109.4]
  reg [63:0] _RAND_11;
  reg [4:0] data_bank; // @[NV_NVDLA_CSC_dl_for_check.scala 172:24:@111.4]
  reg [31:0] _RAND_12;
  reg [13:0] datain_width; // @[NV_NVDLA_CSC_dl_for_check.scala 173:27:@113.4]
  reg [31:0] _RAND_13;
  reg [12:0] datain_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 174:31:@115.4]
  reg [31:0] _RAND_14;
  reg [12:0] datain_height_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 175:32:@117.4]
  reg [31:0] _RAND_15;
  reg [10:0] datain_channel_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 176:33:@119.4]
  reg [31:0] _RAND_16;
  reg [2:0] sub_h_total_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 177:29:@120.4]
  reg [31:0] _RAND_17;
  reg [2:0] sub_h_total_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 178:29:@121.4]
  reg [31:0] _RAND_18;
  reg [2:0] sub_h_total_g3; // @[NV_NVDLA_CSC_dl_for_check.scala 180:29:@123.4]
  reg [31:0] _RAND_19;
  reg [2:0] sub_h_total_g4; // @[NV_NVDLA_CSC_dl_for_check.scala 181:29:@124.4]
  reg [31:0] _RAND_20;
  reg [2:0] sub_h_total_g5; // @[NV_NVDLA_CSC_dl_for_check.scala 182:29:@125.4]
  reg [31:0] _RAND_21;
  reg [2:0] sub_h_total_g6; // @[NV_NVDLA_CSC_dl_for_check.scala 183:29:@126.4]
  reg [31:0] _RAND_22;
  reg [2:0] sub_h_total_g8; // @[NV_NVDLA_CSC_dl_for_check.scala 185:29:@128.4]
  reg [31:0] _RAND_23;
  reg [2:0] sub_h_total_g9; // @[NV_NVDLA_CSC_dl_for_check.scala 186:29:@129.4]
  reg [31:0] _RAND_24;
  reg [2:0] sub_h_total_g11; // @[NV_NVDLA_CSC_dl_for_check.scala 188:30:@131.4]
  reg [31:0] _RAND_25;
  reg [2:0] sub_h_cmp_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 189:27:@132.4]
  reg [31:0] _RAND_26;
  reg [2:0] sub_h_cmp_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 190:27:@133.4]
  reg [31:0] _RAND_27;
  reg [3:0] conv_x_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 191:28:@135.4]
  reg [31:0] _RAND_28;
  reg [3:0] conv_y_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 192:28:@137.4]
  reg [31:0] _RAND_29;
  reg [4:0] batch_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 194:24:@140.4]
  reg [31:0] _RAND_30;
  reg [6:0] pixel_x_init; // @[NV_NVDLA_CSC_dl_for_check.scala 195:27:@142.4]
  reg [31:0] _RAND_31;
  reg [6:0] pixel_x_init_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 196:34:@144.4]
  reg [31:0] _RAND_32;
  reg [7:0] pixel_x_add; // @[NV_NVDLA_CSC_dl_for_check.scala 197:26:@146.4]
  reg [31:0] _RAND_33;
  reg [6:0] pixel_x_byte_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 198:34:@148.4]
  reg [31:0] _RAND_34;
  reg [11:0] pixel_ch_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 199:30:@150.4]
  reg [31:0] _RAND_35;
  reg [5:0] x_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 200:23:@152.4]
  reg [31:0] _RAND_36;
  reg [5:0] y_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 201:23:@154.4]
  reg [31:0] _RAND_37;
  reg [15:0] pad_value; // @[NV_NVDLA_CSC_dl_for_check.scala 202:24:@156.4]
  reg [31:0] _RAND_38;
  reg [14:0] entries_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 203:26:@158.4]
  reg [31:0] _RAND_39;
  reg [14:0] h_bias_2_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 204:30:@160.4]
  reg [31:0] _RAND_40;
  reg [14:0] h_bias_3_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 205:30:@162.4]
  reg [31:0] _RAND_41;
  reg [13:0] last_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 207:26:@164.4]
  reg [31:0] _RAND_42;
  reg [14:0] last_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 208:27:@166.4]
  reg [31:0] _RAND_43;
  wire [33:0] _T_670; // @[Bitwise.scala 72:12:@174.6]
  wire [5:0] _T_672; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@176.6]
  wire [4:0] _T_673; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@177.6]
  wire [13:0] _T_675; // @[NV_NVDLA_CSC_dl_for_check.scala 216:48:@179.6]
  wire [6:0] _T_681; // @[NV_NVDLA_CSC_dl_for_check.scala 219:93:@184.6]
  wire [10:0] _T_682; // @[Cat.scala 30:58:@185.6]
  wire [14:0] _T_686; // @[Cat.scala 30:58:@218.6]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [4:0] _GEN_2; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [13:0] _GEN_3; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [12:0] _GEN_4; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [12:0] _GEN_5; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [10:0] _GEN_6; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_7; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_8; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_10; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_11; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_12; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_13; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_15; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_19; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [2:0] _GEN_20; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [3:0] _GEN_21; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [5:0] _GEN_24; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [6:0] _GEN_26; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [6:0] _GEN_27; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [11:0] _GEN_30; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [5:0] _GEN_31; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [14:0] _GEN_34; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [14:0] _GEN_35; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [14:0] _GEN_36; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [13:0] _GEN_37; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [13:0] _GEN_39; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [12:0] _GEN_40; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  wire [11:0] _GEN_43; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  wire [11:0] _GEN_44; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  wire [14:0] _GEN_45; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  wire [14:0] _GEN_46; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  wire [14:0] _GEN_47; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  wire [13:0] _GEN_48; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@238.4]
  wire [14:0] _GEN_49; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@238.4]
  reg [14:0] dat_entry_st; // @[NV_NVDLA_CSC_dl_for_check.scala 287:59:@250.4]
  reg [31:0] _RAND_44;
  wire  _T_763; // @[NV_NVDLA_CSC_dl_for_check.scala 328:37:@313.4]
  wire  _T_764; // @[NV_NVDLA_CSC_dl_for_check.scala 328:23:@314.4]
  wire  _T_1627; // @[NV_NVDLA_CSC_dl_for_check.scala 918:32:@1216.4]
  reg  dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1184.4]
  reg [31:0] _RAND_45;
  wire  _T_1628; // @[NV_NVDLA_CSC_dl_for_check.scala 918:36:@1217.4]
  wire  _T_1629; // @[NV_NVDLA_CSC_dl_for_check.scala 919:35:@1218.4]
  reg  dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1182.4]
  reg [31:0] _RAND_46;
  wire  _T_1630; // @[NV_NVDLA_CSC_dl_for_check.scala 919:39:@1219.4]
  wire  _T_1631; // @[NV_NVDLA_CSC_dl_for_check.scala 918:57:@1220.4]
  wire  _T_1632; // @[NV_NVDLA_CSC_dl_for_check.scala 920:35:@1221.4]
  reg  dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1181.4]
  reg [31:0] _RAND_47;
  wire  _T_1633; // @[NV_NVDLA_CSC_dl_for_check.scala 920:39:@1222.4]
  wire  dat_rsp_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 919:60:@1223.4]
  wire  _T_1635; // @[NV_NVDLA_CSC_dl_for_check.scala 927:42:@1225.4]
  wire [26:0] _T_1639; // @[Bitwise.scala 72:12:@1227.4]
  reg [26:0] _T_1617; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1189.4]
  reg [31:0] _RAND_48;
  wire [26:0] _T_1640; // @[NV_NVDLA_CSC_dl_for_check.scala 927:47:@1228.4]
  wire  _T_1641; // @[NV_NVDLA_CSC_dl_for_check.scala 928:42:@1229.4]
  wire [26:0] _T_1645; // @[Bitwise.scala 72:12:@1231.4]
  reg [26:0] _T_1611; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1187.4]
  reg [31:0] _RAND_49;
  wire [26:0] _T_1646; // @[NV_NVDLA_CSC_dl_for_check.scala 928:47:@1232.4]
  wire [26:0] _T_1647; // @[NV_NVDLA_CSC_dl_for_check.scala 927:66:@1233.4]
  wire  _T_1648; // @[NV_NVDLA_CSC_dl_for_check.scala 929:42:@1234.4]
  wire [26:0] _T_1652; // @[Bitwise.scala 72:12:@1236.4]
  reg [26:0] _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1186.4]
  reg [31:0] _RAND_50;
  wire [26:0] _T_1653; // @[NV_NVDLA_CSC_dl_for_check.scala 929:47:@1237.4]
  wire [26:0] dat_rsp_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 928:66:@1238.4]
  wire  dat_rsp_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 953:26:@1257.4]
  wire  sub_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 325:29:@312.4]
  wire  _T_766; // @[NV_NVDLA_CSC_dl_for_check.scala 328:66:@315.4]
  wire  _T_767; // @[NV_NVDLA_CSC_dl_for_check.scala 328:53:@316.4]
  wire  dat_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 328:42:@317.4]
  wire [13:0] sc2cdma_dat_slices_w; // @[NV_NVDLA_CSC_dl_for_check.scala 329:28:@319.4]
  wire [14:0] sc2cdma_dat_entries_w; // @[NV_NVDLA_CSC_dl_for_check.scala 330:29:@321.4]
  wire [14:0] dat_entry_avl_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 297:28:@261.4]
  wire [15:0] _T_720; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@268.4]
  wire [14:0] dat_entry_st_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@269.4]
  wire [13:0] _T_726; // @[Cat.scala 30:58:@271.4]
  wire [14:0] _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@272.4]
  wire [15:0] _T_727; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@272.4]
  wire [15:0] _T_728; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@273.4]
  wire [14:0] dat_entry_st_inc_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@274.4]
  wire  is_dat_entry_st_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 304:45:@277.4]
  wire [14:0] _T_736; // @[NV_NVDLA_CSC_dl_for_check.scala 305:83:@278.4]
  wire [14:0] dat_entry_st_w; // @[NV_NVDLA_CSC_dl_for_check.scala 305:25:@279.4]
  wire  _T_758; // @[NV_NVDLA_CSC_dl_for_check.scala 316:13:@302.4]
  wire [14:0] _GEN_52; // @[NV_NVDLA_CSC_dl_for_check.scala 316:25:@303.4]
  reg  _T_773; // @[NV_NVDLA_CSC_dl_for_check.scala 332:31:@323.4]
  reg [31:0] _RAND_51;
  reg [13:0] _T_776; // @[Reg.scala 19:20:@326.4]
  reg [31:0] _RAND_52;
  wire [13:0] _GEN_54; // @[Reg.scala 20:19:@327.4]
  reg [14:0] _T_779; // @[Reg.scala 19:20:@331.4]
  reg [31:0] _RAND_53;
  wire [14:0] _GEN_55; // @[Reg.scala 20:19:@332.4]
  reg  _T_784; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@337.4]
  reg [31:0] _RAND_54;
  reg  _T_787; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@338.4]
  reg [31:0] _RAND_55;
  reg  _T_790; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@339.4]
  reg [31:0] _RAND_56;
  reg  _T_793; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@340.4]
  reg [31:0] _RAND_57;
  reg  dl_in_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 345:50:@341.4]
  reg [31:0] _RAND_58;
  reg  _T_817; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@371.4]
  reg [31:0] _RAND_59;
  reg  _T_820; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@372.4]
  reg [31:0] _RAND_60;
  reg  _T_823; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@373.4]
  reg [31:0] _RAND_61;
  reg  _T_826; // @[NV_NVDLA_CSC_dl_for_check.scala 364:36:@374.4]
  reg [31:0] _RAND_62;
  reg [30:0] _T_831; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@376.4]
  reg [31:0] _RAND_63;
  reg [30:0] _T_834; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@377.4]
  reg [31:0] _RAND_64;
  reg [30:0] _T_837; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@378.4]
  reg [31:0] _RAND_65;
  reg [30:0] _T_840; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@379.4]
  reg [31:0] _RAND_66;
  wire [30:0] _T_828; // @[NV_NVDLA_CSC_dl_for_check.scala 365:19:@375.4 NV_NVDLA_CSC_dl_for_check.scala 369:12:@381.4]
  wire [30:0] _GEN_61; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@383.4]
  wire [30:0] _GEN_62; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@387.4]
  wire [30:0] _GEN_63; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@391.4]
  wire [30:0] _GEN_64; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@395.4]
  wire  _T_841; // @[NV_NVDLA_CSC_dl_for_check.scala 378:30:@398.4]
  wire  _T_842; // @[NV_NVDLA_CSC_dl_for_check.scala 378:34:@399.4]
  wire  _T_843; // @[NV_NVDLA_CSC_dl_for_check.scala 379:30:@400.4]
  wire  _T_844; // @[NV_NVDLA_CSC_dl_for_check.scala 379:34:@401.4]
  wire  _T_845; // @[NV_NVDLA_CSC_dl_for_check.scala 378:50:@402.4]
  wire  _T_846; // @[NV_NVDLA_CSC_dl_for_check.scala 380:30:@403.4]
  wire  _T_847; // @[NV_NVDLA_CSC_dl_for_check.scala 380:34:@404.4]
  wire  dl_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 379:50:@405.4]
  wire  _T_848; // @[NV_NVDLA_CSC_dl_for_check.scala 382:37:@406.4]
  wire [30:0] _T_852; // @[Bitwise.scala 72:12:@408.4]
  wire [30:0] _T_853; // @[NV_NVDLA_CSC_dl_for_check.scala 382:42:@409.4]
  wire  _T_854; // @[NV_NVDLA_CSC_dl_for_check.scala 383:37:@410.4]
  wire [30:0] _T_858; // @[Bitwise.scala 72:12:@412.4]
  wire [30:0] _T_859; // @[NV_NVDLA_CSC_dl_for_check.scala 383:42:@413.4]
  wire [30:0] _T_860; // @[NV_NVDLA_CSC_dl_for_check.scala 382:56:@414.4]
  wire  _T_861; // @[NV_NVDLA_CSC_dl_for_check.scala 384:37:@415.4]
  wire [30:0] _T_865; // @[Bitwise.scala 72:12:@417.4]
  wire [30:0] _T_866; // @[NV_NVDLA_CSC_dl_for_check.scala 384:42:@418.4]
  wire [30:0] dl_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 383:56:@419.4]
  wire [4:0] dl_w_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 387:24:@420.4]
  wire [4:0] dl_h_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 388:24:@421.4]
  wire [6:0] dl_channel_size; // @[NV_NVDLA_CSC_dl_for_check.scala 389:28:@422.4]
  wire [6:0] dl_stripe_length; // @[NV_NVDLA_CSC_dl_for_check.scala 390:29:@423.4]
  wire [1:0] dl_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 391:25:@424.4]
  wire  dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 392:25:@425.4]
  wire  dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 393:27:@426.4]
  wire  dl_group_end; // @[NV_NVDLA_CSC_dl_for_check.scala 394:25:@427.4]
  wire  dl_layer_end; // @[NV_NVDLA_CSC_dl_for_check.scala 395:25:@428.4]
  wire  dl_dat_release; // @[NV_NVDLA_CSC_dl_for_check.scala 396:27:@429.4]
  reg [5:0] batch_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 401:24:@432.4]
  reg [31:0] _RAND_67;
  wire [6:0] _T_874; // @[NV_NVDLA_CSC_dl_for_check.scala 405:24:@433.4]
  wire [5:0] _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 407:27:@438.4]
  wire  is_batch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 407:27:@438.4]
  wire [6:0] _T_875; // @[NV_NVDLA_CSC_dl_for_check.scala 404:17:@434.4]
  wire [6:0] _T_876; // @[NV_NVDLA_CSC_dl_for_check.scala 403:17:@435.4]
  wire [5:0] _T_877; // @[NV_NVDLA_CSC_dl_for_check.scala 405:32:@436.4]
  reg [1:0] sub_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 410:24:@440.4]
  reg [31:0] _RAND_68;
  wire [2:0] sub_h_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 413:31:@442.4]
  wire  is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 414:32:@443.4]
  wire  _T_885; // @[NV_NVDLA_CSC_dl_for_check.scala 415:61:@445.4]
  reg [6:0] stripe_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 421:25:@453.4]
  reg [31:0] _RAND_69;
  wire  _T_921; // @[NV_NVDLA_CSC_dl_for_check.scala 448:37:@482.4]
  wire  _T_922; // @[NV_NVDLA_CSC_dl_for_check.scala 448:24:@483.4]
  wire  _T_924; // @[NV_NVDLA_CSC_dl_for_check.scala 448:56:@484.4]
  wire  _T_925; // @[NV_NVDLA_CSC_dl_for_check.scala 448:44:@485.4]
  wire  _T_926; // @[NV_NVDLA_CSC_dl_for_check.scala 448:42:@486.4]
  wire  _T_928; // @[NV_NVDLA_CSC_dl_for_check.scala 448:75:@487.4]
  wire  _T_929; // @[NV_NVDLA_CSC_dl_for_check.scala 448:63:@488.4]
  wire  _T_930; // @[NV_NVDLA_CSC_dl_for_check.scala 448:61:@489.4]
  reg  dat_exec_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 440:32:@475.4]
  reg [31:0] _RAND_70;
  wire  _T_932; // @[NV_NVDLA_CSC_dl_for_check.scala 448:22:@490.4]
  wire  dat_exec_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 447:22:@491.4]
  wire  _T_886; // @[NV_NVDLA_CSC_dl_for_check.scala 415:66:@446.4]
  wire  sub_h_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 415:33:@447.4]
  wire  _T_887; // @[NV_NVDLA_CSC_dl_for_check.scala 417:31:@449.6]
  wire [2:0] _T_889; // @[NV_NVDLA_CSC_dl_for_check.scala 417:21:@450.6]
  wire [2:0] _GEN_65; // @[NV_NVDLA_CSC_dl_for_check.scala 416:23:@448.4]
  wire [7:0] stripe_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 425:33:@456.4]
  wire [7:0] _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 426:51:@457.4]
  wire  _T_895; // @[NV_NVDLA_CSC_dl_for_check.scala 426:51:@457.4]
  wire  is_stripe_equal; // @[NV_NVDLA_CSC_dl_for_check.scala 426:33:@458.4]
  wire  is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 427:34:@460.4]
  wire  _T_898; // @[NV_NVDLA_CSC_dl_for_check.scala 428:52:@462.4]
  wire  stripe_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 428:34:@463.4]
  wire  _T_900; // @[NV_NVDLA_CSC_dl_for_check.scala 432:41:@465.6]
  wire  _T_901; // @[NV_NVDLA_CSC_dl_for_check.scala 432:39:@466.6]
  wire [7:0] _T_903; // @[NV_NVDLA_CSC_dl_for_check.scala 433:22:@467.6]
  wire [7:0] _T_904; // @[NV_NVDLA_CSC_dl_for_check.scala 432:22:@468.6]
  wire [7:0] _T_905; // @[NV_NVDLA_CSC_dl_for_check.scala 431:22:@469.6]
  wire [7:0] _GEN_66; // @[NV_NVDLA_CSC_dl_for_check.scala 430:24:@464.4]
  reg  dat_pipe_local_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 438:35:@473.4]
  reg [31:0] _RAND_71;
  reg  dat_pipe_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 439:32:@474.4]
  reg [31:0] _RAND_72;
  wire  dat_pipe_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 446:27:@480.4]
  wire  _T_914; // @[NV_NVDLA_CSC_dl_for_check.scala 443:49:@477.4]
  wire  _T_917; // @[NV_NVDLA_CSC_dl_for_check.scala 444:32:@478.4]
  wire  dat_pipe_local_valid_w; // @[NV_NVDLA_CSC_dl_for_check.scala 443:33:@479.4]
  reg [7:0] dat_req_bytes_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 456:31:@496.4]
  reg [31:0] _RAND_73;
  wire [7:0] dat_req_bytes; // @[Cat.scala 30:58:@497.4]
  wire [7:0] _GEN_67; // @[NV_NVDLA_CSC_dl_for_check.scala 458:21:@498.4]
  reg [12:0] dataout_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 464:28:@501.4]
  reg [31:0] _RAND_74;
  reg [12:0] dataout_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 465:28:@502.4]
  reg [31:0] _RAND_75;
  wire [12:0] _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@503.4]
  wire [13:0] _T_941; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@503.4]
  wire [12:0] dataout_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@504.4]
  wire  _T_942; // @[NV_NVDLA_CSC_dl_for_check.scala 469:29:@505.4]
  wire  _T_943; // @[NV_NVDLA_CSC_dl_for_check.scala 469:61:@506.4]
  wire  is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 469:44:@507.4]
  wire  _T_945; // @[NV_NVDLA_CSC_dl_for_check.scala 472:43:@510.4]
  wire  _T_946; // @[NV_NVDLA_CSC_dl_for_check.scala 472:41:@511.4]
  wire [12:0] _T_947; // @[NV_NVDLA_CSC_dl_for_check.scala 473:26:@512.4]
  wire [12:0] _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 472:26:@513.4]
  wire [12:0] dataout_w_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 471:26:@514.4]
  wire  _T_950; // @[NV_NVDLA_CSC_dl_for_check.scala 474:70:@516.4]
  wire  dataout_w_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 474:37:@517.4]
  wire  _T_951; // @[NV_NVDLA_CSC_dl_for_check.scala 475:55:@518.4]
  wire  _T_952; // @[NV_NVDLA_CSC_dl_for_check.scala 475:71:@519.4]
  wire  dataout_w_ori_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 475:37:@520.4]
  wire [12:0] _GEN_68; // @[NV_NVDLA_CSC_dl_for_check.scala 477:27:@521.4]
  wire [12:0] _GEN_69; // @[NV_NVDLA_CSC_dl_for_check.scala 480:27:@524.4]
  reg [10:0] datain_c_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 485:27:@527.4]
  reg [31:0] _RAND_76;
  wire  is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@528.4]
  wire  _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 488:70:@530.4]
  wire  datain_c_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 488:36:@531.4]
  wire [11:0] _T_960; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@533.6]
  wire [10:0] _T_961; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@534.6]
  wire [10:0] _T_962; // @[NV_NVDLA_CSC_dl_for_check.scala 492:24:@535.6]
  wire [10:0] _T_963; // @[NV_NVDLA_CSC_dl_for_check.scala 491:24:@536.6]
  wire [10:0] _GEN_70; // @[NV_NVDLA_CSC_dl_for_check.scala 490:26:@532.4]
  reg [13:0] datain_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 497:27:@539.4]
  reg [31:0] _RAND_77;
  reg [13:0] datain_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 498:27:@540.4]
  reg [31:0] _RAND_78;
  reg [15:0] pixel_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 499:26:@541.4]
  reg [31:0] _RAND_79;
  reg [15:0] pixel_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 500:26:@542.4]
  reg [31:0] _RAND_80;
  reg [15:0] pixel_w_ch_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 501:29:@543.4]
  reg [31:0] _RAND_81;
  reg [12:0] channel_op_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 502:29:@544.4]
  reg [31:0] _RAND_82;
  reg  pixel_force_clr_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 504:33:@546.4]
  reg [31:0] _RAND_83;
  reg  pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 505:35:@547.4]
  reg [31:0] _RAND_84;
  wire [12:0] _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@548.4]
  wire [13:0] _T_983; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@548.4]
  wire [13:0] _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@549.4]
  wire [13:0] datain_w_cnt_st; // @[NV_NVDLA_CSC_dl_for_check.scala 507:26:@550.4]
  wire [13:0] _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@551.4]
  wire [14:0] _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@551.4]
  wire [13:0] datain_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@552.4]
  wire [13:0] _T_988; // @[NV_NVDLA_CSC_dl_for_check.scala 514:25:@555.4]
  wire [13:0] _T_989; // @[NV_NVDLA_CSC_dl_for_check.scala 513:25:@556.4]
  wire [13:0] datain_w_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 512:25:@557.4]
  wire [5:0] _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@558.4]
  wire [10:0] dl_w_offset_ext; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@558.4]
  wire [13:0] _GEN_688; // @[NV_NVDLA_CSC_dl_for_check.scala 517:34:@559.4]
  wire [14:0] _T_990; // @[NV_NVDLA_CSC_dl_for_check.scala 517:34:@559.4]
  wire [13:0] datain_w_cur; // @[NV_NVDLA_CSC_dl_for_check.scala 517:53:@560.4]
  wire  _T_993; // @[NV_NVDLA_CSC_dl_for_check.scala 518:96:@563.4]
  wire  _T_994; // @[NV_NVDLA_CSC_dl_for_check.scala 518:86:@564.4]
  wire  _T_995; // @[NV_NVDLA_CSC_dl_for_check.scala 518:84:@565.4]
  wire  datain_w_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 518:36:@566.4]
  wire  _T_998; // @[NV_NVDLA_CSC_dl_for_check.scala 519:99:@569.4]
  wire  _T_999; // @[NV_NVDLA_CSC_dl_for_check.scala 519:89:@570.4]
  wire  _T_1000; // @[NV_NVDLA_CSC_dl_for_check.scala 519:87:@571.4]
  wire  datain_w_ori_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 519:36:@572.4]
  wire [7:0] pixel_x_cnt_add; // @[NV_NVDLA_CSC_dl_for_check.scala 522:26:@573.4]
  wire  _T_1004; // @[NV_NVDLA_CSC_dl_for_check.scala 524:79:@575.4]
  wire [7:0] _T_1008; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@578.4]
  wire [6:0] _T_1009; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@579.4]
  wire [6:0] total_channel_op; // @[NV_NVDLA_CSC_dl_for_check.scala 524:27:@580.4]
  wire  _T_1010; // @[NV_NVDLA_CSC_dl_for_check.scala 526:37:@581.4]
  wire  _T_1012; // @[NV_NVDLA_CSC_dl_for_check.scala 527:35:@582.4]
  wire [13:0] _T_1014; // @[NV_NVDLA_CSC_dl_for_check.scala 527:66:@583.4]
  wire [13:0] _T_1015; // @[NV_NVDLA_CSC_dl_for_check.scala 527:22:@584.4]
  wire [13:0] _T_1016; // @[NV_NVDLA_CSC_dl_for_check.scala 526:22:@585.4]
  wire [12:0] _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@587.4]
  wire  next_is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@587.4]
  wire  _T_1017; // @[NV_NVDLA_CSC_dl_for_check.scala 533:39:@588.4]
  wire  _T_1018; // @[NV_NVDLA_CSC_dl_for_check.scala 533:54:@589.4]
  wire  _T_1019; // @[NV_NVDLA_CSC_dl_for_check.scala 533:71:@590.4]
  wire  _T_1022; // @[NV_NVDLA_CSC_dl_for_check.scala 534:73:@593.4]
  wire  _T_1023; // @[NV_NVDLA_CSC_dl_for_check.scala 534:71:@594.4]
  wire [15:0] _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@595.4]
  wire [16:0] _T_1024; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@595.4]
  wire  _T_1026; // @[NV_NVDLA_CSC_dl_for_check.scala 535:54:@597.4]
  wire [15:0] _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@598.4]
  wire [16:0] _T_1027; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@598.4]
  wire  _T_1029; // @[NV_NVDLA_CSC_dl_for_check.scala 536:56:@600.4]
  wire  _T_1030; // @[NV_NVDLA_CSC_dl_for_check.scala 536:54:@601.4]
  wire [16:0] _T_1032; // @[NV_NVDLA_CSC_dl_for_check.scala 536:91:@602.4]
  wire  _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 537:41:@603.4]
  wire  _T_1034; // @[NV_NVDLA_CSC_dl_for_check.scala 537:39:@604.4]
  wire [15:0] _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@605.4]
  wire [16:0] _T_1035; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@605.4]
  wire [16:0] _T_1036; // @[NV_NVDLA_CSC_dl_for_check.scala 537:24:@606.4]
  wire [16:0] _T_1037; // @[NV_NVDLA_CSC_dl_for_check.scala 536:24:@607.4]
  wire [16:0] _T_1038; // @[NV_NVDLA_CSC_dl_for_check.scala 535:24:@608.4]
  wire [16:0] _T_1039; // @[NV_NVDLA_CSC_dl_for_check.scala 534:24:@609.4]
  wire [16:0] _T_1040; // @[NV_NVDLA_CSC_dl_for_check.scala 533:24:@610.4]
  wire [16:0] _T_1041; // @[NV_NVDLA_CSC_dl_for_check.scala 532:24:@611.4]
  wire [15:0] pixel_w_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 537:105:@612.4]
  wire [9:0] _T_1047; // @[NV_NVDLA_CSC_dl_for_check.scala 539:68:@614.4]
  wire [14:0] pixel_w_cur; // @[Cat.scala 30:58:@615.4]
  wire  _T_1056; // @[NV_NVDLA_CSC_dl_for_check.scala 542:68:@626.4]
  wire  _T_1057; // @[NV_NVDLA_CSC_dl_for_check.scala 542:57:@627.4]
  wire  _T_1058; // @[NV_NVDLA_CSC_dl_for_check.scala 542:72:@628.4]
  wire  _T_1059; // @[NV_NVDLA_CSC_dl_for_check.scala 542:88:@629.4]
  wire  _T_1060; // @[NV_NVDLA_CSC_dl_for_check.scala 542:103:@630.4]
  wire  pixel_ch_ori_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 542:39:@631.4]
  wire  _T_1062; // @[NV_NVDLA_CSC_dl_for_check.scala 544:42:@633.4]
  wire  _T_1065; // @[NV_NVDLA_CSC_dl_for_check.scala 544:74:@634.4]
  wire  pixel_force_fetch; // @[NV_NVDLA_CSC_dl_for_check.scala 544:28:@635.4]
  wire  _T_1067; // @[NV_NVDLA_CSC_dl_for_check.scala 545:36:@637.4]
  wire  _T_1068; // @[NV_NVDLA_CSC_dl_for_check.scala 545:72:@638.4]
  wire  pixel_force_clr; // @[NV_NVDLA_CSC_dl_for_check.scala 545:51:@639.4]
  wire [13:0] _GEN_71; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@640.4]
  wire [15:0] _GEN_72; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@640.4]
  wire [13:0] _GEN_73; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@644.4]
  wire [15:0] _GEN_74; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@644.4]
  wire [15:0] _GEN_75; // @[NV_NVDLA_CSC_dl_for_check.scala 555:26:@648.4]
  reg [13:0] datain_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 561:27:@651.4]
  reg [31:0] _RAND_85;
  reg [13:0] datain_h_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 562:27:@652.4]
  reg [31:0] _RAND_86;
  wire [13:0] _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@653.4]
  wire [14:0] _T_1074; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@653.4]
  wire [14:0] _T_1075; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@654.4]
  wire [13:0] datain_h_cnt_st; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@655.4]
  wire [13:0] _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@656.4]
  wire [14:0] _T_1076; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@656.4]
  wire [13:0] datain_h_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@657.4]
  wire  _T_1077; // @[NV_NVDLA_CSC_dl_for_check.scala 566:52:@658.4]
  wire  _T_1078; // @[NV_NVDLA_CSC_dl_for_check.scala 566:35:@659.4]
  wire [13:0] _T_1081; // @[NV_NVDLA_CSC_dl_for_check.scala 568:25:@662.4]
  wire [13:0] _T_1082; // @[NV_NVDLA_CSC_dl_for_check.scala 567:25:@663.4]
  wire [13:0] datain_h_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 566:25:@664.4]
  wire  _T_1085; // @[NV_NVDLA_CSC_dl_for_check.scala 569:91:@667.4]
  wire  _T_1086; // @[NV_NVDLA_CSC_dl_for_check.scala 569:54:@668.4]
  wire  datain_h_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 569:36:@669.4]
  wire [5:0] _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@673.4]
  wire [10:0] dl_h_offset_ext; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@673.4]
  wire [13:0] _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 572:34:@674.4]
  wire [14:0] _T_1089; // @[NV_NVDLA_CSC_dl_for_check.scala 572:34:@674.4]
  wire [14:0] _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 572:53:@675.4]
  wire [15:0] _T_1090; // @[NV_NVDLA_CSC_dl_for_check.scala 572:53:@675.4]
  wire [13:0] datain_h_cur; // @[NV_NVDLA_CSC_dl_for_check.scala 572:66:@676.4]
  wire [13:0] _GEN_76; // @[NV_NVDLA_CSC_dl_for_check.scala 574:26:@677.4]
  wire [13:0] _GEN_77; // @[NV_NVDLA_CSC_dl_for_check.scala 575:26:@680.4]
  wire  _T_1091; // @[NV_NVDLA_CSC_dl_for_check.scala 578:39:@683.4]
  wire [13:0] _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@684.4]
  wire  _T_1092; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@684.4]
  wire  _T_1093; // @[NV_NVDLA_CSC_dl_for_check.scala 578:44:@685.4]
  wire  _T_1094; // @[NV_NVDLA_CSC_dl_for_check.scala 578:92:@686.4]
  wire  _T_1095; // @[NV_NVDLA_CSC_dl_for_check.scala 578:78:@687.4]
  wire [13:0] _GEN_699; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@688.4]
  wire  _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@688.4]
  wire  dat_conv_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 578:97:@689.4]
  wire  dat_img_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 581:42:@699.4]
  wire  _T_1179; // @[NV_NVDLA_CSC_dl_for_check.scala 666:33:@785.4]
  wire  _T_1180; // @[NV_NVDLA_CSC_dl_for_check.scala 667:24:@786.4]
  wire [12:0] _T_1182; // @[NV_NVDLA_CSC_dl_for_check.scala 667:77:@787.4]
  wire [14:0] _T_1183; // @[Cat.scala 30:58:@788.4]
  wire  _T_1185; // @[NV_NVDLA_CSC_dl_for_check.scala 668:38:@789.4]
  wire [11:0] _T_1190; // @[NV_NVDLA_CSC_dl_for_check.scala 669:54:@792.4]
  wire [14:0] _T_1191; // @[Cat.scala 30:58:@793.4]
  wire [14:0] _T_1192; // @[NV_NVDLA_CSC_dl_for_check.scala 668:23:@794.4]
  wire [14:0] _T_1193; // @[NV_NVDLA_CSC_dl_for_check.scala 667:23:@795.4]
  wire [14:0] w_bias_int8; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@796.4]
  wire [13:0] w_bias_w; // @[NV_NVDLA_CSC_dl_for_check.scala 678:24:@798.4]
  wire [11:0] _T_1108; // @[NV_NVDLA_CSC_dl_for_check.scala 585:32:@701.4]
  wire [14:0] _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@702.4]
  wire  dat_img_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@702.4]
  wire  _T_1109; // @[NV_NVDLA_CSC_dl_for_check.scala 586:34:@703.4]
  wire  dat_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 586:24:@704.4]
  wire  _T_1110; // @[NV_NVDLA_CSC_dl_for_check.scala 587:29:@705.4]
  wire  dat_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 587:33:@706.4]
  wire  _T_1111; // @[NV_NVDLA_CSC_dl_for_check.scala 588:39:@707.4]
  wire  _T_1112; // @[NV_NVDLA_CSC_dl_for_check.scala 588:37:@708.4]
  wire  _T_1113; // @[NV_NVDLA_CSC_dl_for_check.scala 588:56:@709.4]
  wire  dat_req_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 588:54:@710.4]
  wire  _T_1114; // @[NV_NVDLA_CSC_dl_for_check.scala 591:37:@711.4]
  wire  _T_1115; // @[NV_NVDLA_CSC_dl_for_check.scala 591:27:@712.4]
  wire  _T_1116; // @[NV_NVDLA_CSC_dl_for_check.scala 591:54:@713.4]
  wire  dat_req_sub_c_w; // @[NV_NVDLA_CSC_dl_for_check.scala 591:26:@714.4]
  wire [1:0] dat_req_sub_w_w; // @[NV_NVDLA_CSC_dl_for_check.scala 592:35:@715.4]
  wire  _T_1118; // @[NV_NVDLA_CSC_dl_for_check.scala 593:55:@716.4]
  wire  dat_req_sub_w_st_en; // @[NV_NVDLA_CSC_dl_for_check.scala 593:42:@717.4]
  wire  dat_req_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 596:42:@719.4]
  wire [9:0] dat_req_flag_w; // @[Cat.scala 30:58:@723.4]
  reg  dat_req_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 603:31:@724.4]
  reg [31:0] _RAND_87;
  reg [1:0] dat_req_sub_w_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 604:31:@725.4]
  reg [31:0] _RAND_88;
  reg [1:0] dat_req_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 605:31:@726.4]
  reg [31:0] _RAND_89;
  reg  dat_req_sub_c_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 606:31:@727.4]
  reg [31:0] _RAND_90;
  reg  dat_req_ch_end_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:32:@728.4]
  reg [31:0] _RAND_91;
  reg  dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 608:31:@729.4]
  reg [31:0] _RAND_92;
  reg [1:0] dat_req_cur_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 609:35:@730.4]
  reg [31:0] _RAND_93;
  reg  dat_req_sub_w_st_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 610:34:@731.4]
  reg [31:0] _RAND_94;
  reg [8:0] dat_req_flag_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 611:30:@732.4]
  reg [31:0] _RAND_95;
  reg  dat_req_rls_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 612:29:@733.4]
  reg [31:0] _RAND_96;
  wire  _T_1142; // @[NV_NVDLA_CSC_dl_for_check.scala 623:38:@743.6]
  wire  _T_1143; // @[NV_NVDLA_CSC_dl_for_check.scala 623:56:@744.6]
  wire [1:0] _GEN_78; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire [1:0] _GEN_79; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_80; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_81; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_82; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire [1:0] _GEN_83; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire [9:0] _GEN_84; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_85; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_86; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_87; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  wire  _GEN_88; // @[NV_NVDLA_CSC_dl_for_check.scala 627:26:@749.4]
  reg [12:0] c_bias; // @[NV_NVDLA_CSC_dl_for_check.scala 635:21:@752.4]
  reg [31:0] _RAND_97;
  reg [12:0] c_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 636:24:@753.4]
  reg [31:0] _RAND_98;
  reg [12:0] h_bias_0_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 637:26:@754.4]
  reg [31:0] _RAND_99;
  reg [12:0] h_bias_1_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 638:26:@755.4]
  reg [31:0] _RAND_100;
  reg [12:0] h_bias_2_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 639:26:@756.4]
  reg [31:0] _RAND_101;
  reg [12:0] h_bias_3_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 640:26:@757.4]
  reg [31:0] _RAND_102;
  reg [12:0] w_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 641:24:@758.4]
  reg [31:0] _RAND_103;
  wire  _T_1158; // @[NV_NVDLA_CSC_dl_for_check.scala 644:32:@759.4]
  wire  _T_1159; // @[NV_NVDLA_CSC_dl_for_check.scala 644:22:@760.4]
  wire [11:0] _T_1160; // @[NV_NVDLA_CSC_dl_for_check.scala 644:49:@761.4]
  wire [11:0] c_bias_add; // @[NV_NVDLA_CSC_dl_for_check.scala 644:21:@762.4]
  wire  _T_1163; // @[NV_NVDLA_CSC_dl_for_check.scala 646:34:@763.4]
  wire [12:0] _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@764.4]
  wire [13:0] _T_1165; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@764.4]
  wire [12:0] _T_1166; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@765.4]
  wire [12:0] _T_1167; // @[NV_NVDLA_CSC_dl_for_check.scala 646:19:@766.4]
  wire [12:0] c_bias_w; // @[NV_NVDLA_CSC_dl_for_check.scala 645:19:@767.4]
  wire  c_bias_d1_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 648:31:@771.4]
  wire [13:0] _GEN_703; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@772.4]
  wire [25:0] _T_1170; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@772.4]
  wire [12:0] h_bias_0_w; // @[NV_NVDLA_CSC_dl_for_check.scala 651:50:@773.4]
  wire [11:0] _GEN_704; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@774.4]
  wire [16:0] _T_1171; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@774.4]
  wire [12:0] h_bias_1_w; // @[NV_NVDLA_CSC_dl_for_check.scala 652:49:@775.4]
  wire [14:0] _GEN_705; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@776.4]
  wire [20:0] _T_1172; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@776.4]
  wire [12:0] h_bias_2_w; // @[NV_NVDLA_CSC_dl_for_check.scala 653:47:@777.4]
  wire [16:0] _T_1174; // @[NV_NVDLA_CSC_dl_for_check.scala 654:79:@778.4]
  wire [16:0] _T_1175; // @[NV_NVDLA_CSC_dl_for_check.scala 654:21:@779.4]
  wire [12:0] h_bias_3_w; // @[NV_NVDLA_CSC_dl_for_check.scala 654:97:@780.4]
  wire  _T_1176; // @[NV_NVDLA_CSC_dl_for_check.scala 655:45:@781.4]
  wire  _T_1177; // @[NV_NVDLA_CSC_dl_for_check.scala 655:34:@782.4]
  wire [1:0] h_bias_reg_en; // @[Cat.scala 30:58:@783.4]
  wire [12:0] _GEN_89; // @[NV_NVDLA_CSC_dl_for_check.scala 682:20:@800.4]
  wire [12:0] _GEN_90; // @[NV_NVDLA_CSC_dl_for_check.scala 685:23:@803.4]
  wire  _T_1196; // @[NV_NVDLA_CSC_dl_for_check.scala 688:19:@806.4]
  wire [12:0] _GEN_91; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@807.4]
  wire [12:0] _GEN_92; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@807.4]
  wire [12:0] _GEN_93; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@807.4]
  wire  _T_1197; // @[NV_NVDLA_CSC_dl_for_check.scala 693:19:@812.4]
  wire [12:0] _GEN_94; // @[NV_NVDLA_CSC_dl_for_check.scala 693:23:@813.4]
  wire [13:0] _GEN_95; // @[NV_NVDLA_CSC_dl_for_check.scala 696:20:@816.4]
  reg [12:0] dat_req_sub_h_addr_0; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@828.4]
  reg [31:0] _RAND_104;
  reg [12:0] dat_req_sub_h_addr_1; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@828.4]
  reg [31:0] _RAND_105;
  reg [12:0] dat_req_sub_h_addr_2; // @[NV_NVDLA_CSC_dl_for_check.scala 704:33:@828.4]
  reg [31:0] _RAND_106;
  reg  sc2buf_dat_rd_en_out; // @[NV_NVDLA_CSC_dl_for_check.scala 705:35:@829.4]
  reg [31:0] _RAND_107;
  reg [17:0] sc2buf_dat_rd_addr_out; // @[NV_NVDLA_CSC_dl_for_check.scala 706:37:@831.4]
  reg [31:0] _RAND_108;
  reg  dat_req_pipe_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 707:32:@832.4]
  reg [31:0] _RAND_109;
  reg [1:0] dat_req_pipe_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 709:33:@834.4]
  reg [31:0] _RAND_110;
  reg [1:0] dat_req_pipe_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 710:33:@835.4]
  reg [31:0] _RAND_111;
  reg  dat_req_pipe_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 711:33:@836.4]
  reg [31:0] _RAND_112;
  reg  dat_req_pipe_ch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 712:34:@837.4]
  reg [31:0] _RAND_113;
  reg [7:0] dat_req_pipe_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 713:33:@838.4]
  reg [31:0] _RAND_114;
  reg  dat_req_pipe_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 714:33:@839.4]
  reg [31:0] _RAND_115;
  reg [1:0] dat_req_pipe_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 715:37:@840.4]
  reg [31:0] _RAND_116;
  reg  dat_req_pipe_sub_w_st; // @[NV_NVDLA_CSC_dl_for_check.scala 716:36:@841.4]
  reg [31:0] _RAND_117;
  reg  dat_req_pipe_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 717:31:@842.4]
  reg [31:0] _RAND_118;
  reg [8:0] dat_req_pipe_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 718:32:@843.4]
  reg [31:0] _RAND_119;
  wire [13:0] _T_1288; // @[NV_NVDLA_CSC_dl_for_check.scala 720:30:@844.4]
  wire [13:0] _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 720:45:@845.4]
  wire [14:0] _T_1289; // @[NV_NVDLA_CSC_dl_for_check.scala 720:45:@845.4]
  wire [14:0] _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 720:60:@846.4]
  wire [15:0] _T_1290; // @[NV_NVDLA_CSC_dl_for_check.scala 720:60:@846.4]
  wire [12:0] h_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 720:75:@847.4]
  wire [14:0] _GEN_709; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@848.4]
  wire [15:0] _T_1291; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@848.4]
  wire [15:0] _GEN_710; // @[NV_NVDLA_CSC_dl_for_check.scala 721:53:@849.4]
  wire [16:0] _T_1292; // @[NV_NVDLA_CSC_dl_for_check.scala 721:53:@849.4]
  wire [16:0] _GEN_711; // @[NV_NVDLA_CSC_dl_for_check.scala 721:66:@850.4]
  wire [17:0] dat_req_addr_sum; // @[NV_NVDLA_CSC_dl_for_check.scala 721:66:@850.4]
  wire [17:0] _GEN_712; // @[NV_NVDLA_CSC_dl_for_check.scala 722:45:@853.4]
  wire  is_dat_req_addr_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 722:45:@853.4]
  wire [18:0] _T_1305; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@856.4]
  wire [18:0] _T_1306; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@857.4]
  wire [17:0] dat_req_addr_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@858.4]
  wire  _T_1307; // @[NV_NVDLA_CSC_dl_for_check.scala 724:35:@859.4]
  wire [12:0] _T_1313; // @[NV_NVDLA_CSC_dl_for_check.scala 725:83:@861.4]
  wire [17:0] _T_1314; // @[NV_NVDLA_CSC_dl_for_check.scala 725:25:@862.4]
  wire [17:0] dat_req_addr_w; // @[NV_NVDLA_CSC_dl_for_check.scala 724:25:@863.4]
  wire  _T_1333; // @[Mux.scala 46:19:@873.4]
  wire [12:0] _T_1334; // @[Mux.scala 46:16:@874.4]
  wire  _T_1335; // @[Mux.scala 46:19:@875.4]
  wire [12:0] _T_1336; // @[Mux.scala 46:16:@876.4]
  wire  _T_1337; // @[Mux.scala 46:19:@877.4]
  wire [12:0] dat_req_addr_last; // @[Mux.scala 46:16:@878.4]
  wire [17:0] _GEN_715; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@879.4]
  wire  _T_1338; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@879.4]
  wire  _T_1339; // @[NV_NVDLA_CSC_dl_for_check.scala 732:85:@880.4]
  wire  sc2buf_dat_rd_en_w; // @[NV_NVDLA_CSC_dl_for_check.scala 732:43:@881.4]
  wire  _T_1340; // @[NV_NVDLA_CSC_dl_for_check.scala 734:38:@882.4]
  wire  _T_1342; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@883.4]
  wire  _T_1343; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@884.4]
  wire  dat_req_sub_h_addr_en_0; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@885.4]
  wire  _T_1347; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@887.4]
  wire  _T_1348; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@888.4]
  wire  dat_req_sub_h_addr_en_1; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@889.4]
  wire  _T_1352; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@891.4]
  wire  _T_1353; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@892.4]
  wire  dat_req_sub_h_addr_en_2; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@893.4]
  wire [17:0] _GEN_96; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@903.4]
  wire [17:0] _GEN_97; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@906.4]
  wire [17:0] _GEN_98; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@909.4]
  wire  _T_1369; // @[NV_NVDLA_CSC_dl_for_check.scala 747:14:@916.4]
  wire [17:0] _GEN_100; // @[NV_NVDLA_CSC_dl_for_check.scala 747:34:@917.4]
  wire [1:0] _GEN_101; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire [1:0] _GEN_102; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire  _GEN_103; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire  _GEN_104; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire [7:0] _GEN_105; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire  _GEN_106; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire [1:0] _GEN_107; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire  _GEN_108; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire  _GEN_109; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire [8:0] _GEN_110; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  wire [6:0] _T_1379; // @[Cat.scala 30:58:@944.4]
  wire [28:0] dat_req_pipe_pd; // @[Cat.scala 30:58:@950.4]
  reg  _T_1389; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@952.4]
  reg [31:0] _RAND_120;
  reg  _T_1392; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@953.4]
  reg [31:0] _RAND_121;
  reg  _T_1395; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@954.4]
  reg [31:0] _RAND_122;
  reg  _T_1398; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@955.4]
  reg [31:0] _RAND_123;
  reg  _T_1401; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@956.4]
  reg [31:0] _RAND_124;
  reg  dat_rsp_pipe_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 781:73:@957.4]
  reg [31:0] _RAND_125;
  reg [28:0] _T_1408; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@959.4]
  reg [31:0] _RAND_126;
  reg [28:0] _T_1411; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@960.4]
  reg [31:0] _RAND_127;
  reg [28:0] _T_1414; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@961.4]
  reg [31:0] _RAND_128;
  reg [28:0] _T_1417; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@962.4]
  reg [31:0] _RAND_129;
  reg [28:0] _T_1420; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@963.4]
  reg [31:0] _RAND_130;
  reg [28:0] dat_rsp_pipe_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 783:71:@964.4]
  reg [31:0] _RAND_131;
  wire [28:0] _GEN_111; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@992.4]
  wire [28:0] _GEN_114; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1001.4]
  wire [28:0] _GEN_117; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1010.4]
  wire [28:0] _GEN_120; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1019.4]
  wire [28:0] _GEN_123; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1028.4]
  wire [28:0] _GEN_126; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1037.4]
  wire [1:0] dat_rsp_pipe_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 816:41:@1045.4]
  wire [1:0] dat_rsp_pipe_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 817:41:@1046.4]
  wire  dat_rsp_pipe_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 818:41:@1047.4]
  wire  dat_rsp_pipe_ch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 819:42:@1048.4]
  wire [7:0] dat_rsp_pipe_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 820:41:@1049.4]
  wire [1:0] dat_rsp_pipe_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 821:45:@1050.4]
  wire  dat_rsp_pipe_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 824:39:@1053.4]
  wire [8:0] dat_rsp_pipe_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 825:40:@1054.4]
  reg  dat_l0c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 830:29:@1055.4]
  reg [31:0] _RAND_132;
  reg  dat_l0c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 834:29:@1059.4]
  reg [31:0] _RAND_133;
  reg [511:0] dat_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 839:19:@1063.4]
  reg [511:0] _RAND_134;
  reg [511:0] dat_l0c1; // @[NV_NVDLA_CSC_dl_for_check.scala 843:19:@1067.4]
  reg [511:0] _RAND_135;
  wire  _T_1515; // @[NV_NVDLA_CSC_dl_for_check.scala 855:69:@1082.4]
  wire  _T_1516; // @[NV_NVDLA_CSC_dl_for_check.scala 855:74:@1083.4]
  wire  _T_1517; // @[NV_NVDLA_CSC_dl_for_check.scala 855:90:@1084.4]
  wire  dat_l0c1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 855:88:@1085.4]
  wire  _T_1546; // @[NV_NVDLA_CSC_dl_for_check.scala 870:22:@1119.4]
  wire  _T_1560; // @[NV_NVDLA_CSC_dl_for_check.scala 874:48:@1130.4]
  wire  _T_1561; // @[NV_NVDLA_CSC_dl_for_check.scala 874:22:@1131.4]
  reg [7:0] rsp_sft_cnt_l0; // @[NV_NVDLA_CSC_dl_for_check.scala 891:29:@1172.4]
  reg [31:0] _RAND_136;
  reg [7:0] rsp_sft_cnt_l1; // @[NV_NVDLA_CSC_dl_for_check.scala 892:29:@1173.4]
  reg [31:0] _RAND_137;
  reg [7:0] rsp_sft_cnt_l2; // @[NV_NVDLA_CSC_dl_for_check.scala 893:29:@1174.4]
  reg [31:0] _RAND_138;
  reg [7:0] rsp_sft_cnt_l3; // @[NV_NVDLA_CSC_dl_for_check.scala 894:29:@1175.4]
  reg [31:0] _RAND_139;
  reg [7:0] rsp_sft_cnt_l0_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 895:33:@1176.4]
  reg [31:0] _RAND_140;
  reg [7:0] rsp_sft_cnt_l1_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 896:33:@1177.4]
  reg [31:0] _RAND_141;
  reg [7:0] rsp_sft_cnt_l2_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 897:33:@1178.4]
  reg [31:0] _RAND_142;
  reg [7:0] rsp_sft_cnt_l3_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 898:33:@1179.4]
  reg [31:0] _RAND_143;
  reg  dat_rsp_l2_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 903:41:@1183.4]
  reg [31:0] _RAND_144;
  reg [26:0] _T_1614; // @[NV_NVDLA_CSC_dl_for_check.scala 905:41:@1188.4]
  reg [31:0] _RAND_145;
  wire [26:0] _T_1626; // @[Cat.scala 30:58:@1198.4]
  wire [26:0] _GEN_137; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1201.4]
  wire [26:0] _GEN_138; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1205.4]
  wire [26:0] _GEN_139; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1209.4]
  wire [26:0] _GEN_140; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1213.4]
  wire  dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 931:39:@1239.4]
  wire  dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 932:39:@1240.4]
  wire  dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 933:39:@1241.4]
  wire  dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 934:39:@1242.4]
  wire [8:0] dat_rsp_l0_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 936:38:@1243.4]
  wire [8:0] dat_rsp_l1_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 937:38:@1244.4]
  wire [8:0] dat_rsp_l2_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 938:38:@1245.4]
  wire [8:0] dat_rsp_l3_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 939:38:@1246.4]
  wire  dat_rsp_l0_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 941:44:@1247.4]
  wire  dat_rsp_l1_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 942:44:@1248.4]
  wire  dat_rsp_l2_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 943:44:@1249.4]
  wire  dat_rsp_l3_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 944:44:@1250.4]
  wire [1:0] dat_rsp_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 947:31:@1251.4]
  wire [7:0] dat_rsp_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 951:31:@1255.4]
  wire [1:0] dat_rsp_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 952:35:@1256.4]
  wire [8:0] dat_rsp_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 954:30:@1259.4]
  wire [7:0] rsp_sft_cnt_l0_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 963:29:@1265.4]
  wire  _T_1664; // @[NV_NVDLA_CSC_dl_for_check.scala 968:50:@1269.4]
  wire [7:0] _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1270.4]
  wire [8:0] _T_1666; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1270.4]
  wire [8:0] _GEN_717; // @[NV_NVDLA_CSC_dl_for_check.scala 968:134:@1271.4]
  wire [9:0] _T_1667; // @[NV_NVDLA_CSC_dl_for_check.scala 968:134:@1271.4]
  wire [9:0] _T_1668; // @[NV_NVDLA_CSC_dl_for_check.scala 968:134:@1272.4]
  wire [9:0] _T_1669; // @[NV_NVDLA_CSC_dl_for_check.scala 968:29:@1273.4]
  wire [7:0] rsp_sft_cnt_l0_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 968:156:@1274.4]
  wire [8:0] _T_1673; // @[NV_NVDLA_CSC_dl_for_check.scala 969:111:@1276.4]
  wire [9:0] _T_1674; // @[NV_NVDLA_CSC_dl_for_check.scala 969:134:@1277.4]
  wire [9:0] _T_1675; // @[NV_NVDLA_CSC_dl_for_check.scala 969:134:@1278.4]
  wire [9:0] _T_1676; // @[NV_NVDLA_CSC_dl_for_check.scala 969:29:@1279.4]
  wire [7:0] rsp_sft_cnt_l1_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 969:156:@1280.4]
  wire [8:0] _T_1680; // @[NV_NVDLA_CSC_dl_for_check.scala 970:111:@1282.4]
  wire [9:0] _T_1681; // @[NV_NVDLA_CSC_dl_for_check.scala 970:134:@1283.4]
  wire [9:0] _T_1682; // @[NV_NVDLA_CSC_dl_for_check.scala 970:29:@1284.4]
  wire [7:0] rsp_sft_cnt_l2_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 970:156:@1285.4]
  wire [8:0] _T_1686; // @[NV_NVDLA_CSC_dl_for_check.scala 971:111:@1287.4]
  wire [9:0] _T_1687; // @[NV_NVDLA_CSC_dl_for_check.scala 971:134:@1288.4]
  wire [9:0] _T_1688; // @[NV_NVDLA_CSC_dl_for_check.scala 971:29:@1289.4]
  wire [7:0] rsp_sft_cnt_l3_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 971:156:@1290.4]
  wire  _T_1690; // @[NV_NVDLA_CSC_dl_for_check.scala 980:52:@1291.4]
  wire  _T_1691; // @[NV_NVDLA_CSC_dl_for_check.scala 980:50:@1292.4]
  wire  _T_1692; // @[NV_NVDLA_CSC_dl_for_check.scala 981:50:@1293.4]
  wire [7:0] _T_1697; // @[NV_NVDLA_CSC_dl_for_check.scala 981:27:@1296.4]
  wire [7:0] _T_1698; // @[NV_NVDLA_CSC_dl_for_check.scala 980:27:@1297.4]
  wire [7:0] rsp_sft_cnt_l0_w; // @[NV_NVDLA_CSC_dl_for_check.scala 979:27:@1298.4]
  wire  _T_1700; // @[NV_NVDLA_CSC_dl_for_check.scala 985:52:@1299.4]
  wire  _T_1701; // @[NV_NVDLA_CSC_dl_for_check.scala 985:50:@1300.4]
  wire  _T_1702; // @[NV_NVDLA_CSC_dl_for_check.scala 986:50:@1301.4]
  wire [7:0] _T_1707; // @[NV_NVDLA_CSC_dl_for_check.scala 986:27:@1304.4]
  wire [7:0] _T_1708; // @[NV_NVDLA_CSC_dl_for_check.scala 985:27:@1305.4]
  wire [7:0] rsp_sft_cnt_l1_w; // @[NV_NVDLA_CSC_dl_for_check.scala 984:27:@1306.4]
  wire  _T_1710; // @[NV_NVDLA_CSC_dl_for_check.scala 990:52:@1307.4]
  wire  _T_1711; // @[NV_NVDLA_CSC_dl_for_check.scala 990:50:@1308.4]
  wire  _T_1712; // @[NV_NVDLA_CSC_dl_for_check.scala 991:50:@1309.4]
  wire [7:0] _T_1717; // @[NV_NVDLA_CSC_dl_for_check.scala 991:27:@1312.4]
  wire [7:0] _T_1718; // @[NV_NVDLA_CSC_dl_for_check.scala 990:27:@1313.4]
  wire [7:0] rsp_sft_cnt_l2_w; // @[NV_NVDLA_CSC_dl_for_check.scala 989:27:@1314.4]
  wire  _T_1720; // @[NV_NVDLA_CSC_dl_for_check.scala 995:52:@1315.4]
  wire  _T_1721; // @[NV_NVDLA_CSC_dl_for_check.scala 995:50:@1316.4]
  wire  _T_1722; // @[NV_NVDLA_CSC_dl_for_check.scala 996:50:@1317.4]
  wire [7:0] _T_1727; // @[NV_NVDLA_CSC_dl_for_check.scala 996:27:@1320.4]
  wire [7:0] _T_1728; // @[NV_NVDLA_CSC_dl_for_check.scala 995:27:@1321.4]
  wire [7:0] rsp_sft_cnt_l3_w; // @[NV_NVDLA_CSC_dl_for_check.scala 994:27:@1322.4]
  wire  _T_1729; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:46:@1323.4]
  wire  _T_1730; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:51:@1324.4]
  wire  rsp_sft_cnt_l0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:34:@1325.4]
  wire  _T_1731; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:46:@1326.4]
  wire  _T_1732; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:51:@1327.4]
  wire  _T_1734; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:87:@1328.4]
  wire  _T_1735; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:69:@1329.4]
  wire  rsp_sft_cnt_l1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:34:@1330.4]
  wire  _T_1736; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:46:@1331.4]
  wire  _T_1737; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:51:@1332.4]
  wire  _T_1739; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:87:@1333.4]
  wire  _T_1740; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:69:@1334.4]
  wire  rsp_sft_cnt_l2_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:34:@1335.4]
  wire  _T_1741; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:46:@1336.4]
  wire  _T_1742; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:51:@1337.4]
  wire  _T_1745; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:69:@1339.4]
  wire  rsp_sft_cnt_l3_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:34:@1340.4]
  wire  _T_1746; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:50:@1341.4]
  wire  _T_1747; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:55:@1342.4]
  wire  _T_1748; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:73:@1343.4]
  wire  _T_1749; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:97:@1344.4]
  wire  rsp_sft_cnt_l0_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:38:@1345.4]
  wire  _T_1750; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:50:@1346.4]
  wire  _T_1751; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:55:@1347.4]
  wire  _T_1752; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:73:@1348.4]
  wire  _T_1753; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:97:@1349.4]
  wire  _T_1755; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:138:@1350.4]
  wire  _T_1756; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:120:@1351.4]
  wire  rsp_sft_cnt_l1_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:38:@1352.4]
  wire  _T_1757; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:50:@1353.4]
  wire  _T_1758; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:55:@1354.4]
  wire  _T_1759; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:73:@1355.4]
  wire  _T_1760; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:97:@1356.4]
  wire  _T_1762; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:138:@1357.4]
  wire  _T_1763; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:120:@1358.4]
  wire  rsp_sft_cnt_l2_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:38:@1359.4]
  wire  _T_1764; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:50:@1360.4]
  wire  _T_1765; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:55:@1361.4]
  wire  _T_1766; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:73:@1362.4]
  wire  _T_1767; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:97:@1363.4]
  wire  _T_1770; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:120:@1365.4]
  wire  rsp_sft_cnt_l3_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:38:@1366.4]
  wire [7:0] _GEN_141; // @[NV_NVDLA_CSC_dl_for_check.scala 1010:24:@1367.4]
  wire [7:0] _GEN_142; // @[NV_NVDLA_CSC_dl_for_check.scala 1011:24:@1370.4]
  wire [7:0] _GEN_143; // @[NV_NVDLA_CSC_dl_for_check.scala 1012:24:@1373.4]
  wire [7:0] _GEN_144; // @[NV_NVDLA_CSC_dl_for_check.scala 1013:24:@1376.4]
  wire [7:0] _GEN_145; // @[NV_NVDLA_CSC_dl_for_check.scala 1014:28:@1379.4]
  wire [7:0] _GEN_146; // @[NV_NVDLA_CSC_dl_for_check.scala 1015:28:@1382.4]
  wire [7:0] _GEN_147; // @[NV_NVDLA_CSC_dl_for_check.scala 1016:28:@1385.4]
  wire [7:0] _GEN_148; // @[NV_NVDLA_CSC_dl_for_check.scala 1017:28:@1388.4]
  wire [7:0] _T_1771; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:55:@1391.4]
  wire [63:0] _T_1774; // @[Cat.scala 30:58:@1394.4]
  wire [127:0] _T_1775; // @[Cat.scala 30:58:@1395.4]
  wire [255:0] _T_1776; // @[Cat.scala 30:58:@1396.4]
  wire [511:0] dat_rsp_pad_value; // @[Cat.scala 30:58:@1397.4]
  wire [511:0] dat_rsp_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1028:23:@1398.4]
  wire [511:0] dat_rsp_l0c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1033:23:@1402.4]
  wire  _T_1778; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:37:@1407.4]
  wire  _T_1781; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:43:@1408.4]
  wire  _T_1782; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:87:@1409.4]
  wire  _T_1784; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:91:@1410.4]
  wire  _T_1785; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:72:@1411.4]
  wire [255:0] _T_1787; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:171:@1412.4]
  wire [511:0] _T_1788; // @[Cat.scala 30:58:@1413.4]
  wire  _T_1794; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:72:@1417.4]
  wire [255:0] _T_1796; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:171:@1418.4]
  wire [511:0] _T_1797; // @[Cat.scala 30:58:@1419.4]
  wire [511:0] _T_1798; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:27:@1420.4]
  wire [511:0] _T_1799; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:27:@1421.4]
  wire [511:0] dat_rsp_conv_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:27:@1422.4]
  wire [7:0] dat_rsp_conv_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1425.4]
  wire [7:0] dat_rsp_conv_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1427.4]
  wire [7:0] dat_rsp_conv_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1429.4]
  wire [7:0] dat_rsp_conv_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1431.4]
  wire [7:0] dat_rsp_conv_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1433.4]
  wire [7:0] dat_rsp_conv_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1435.4]
  wire [7:0] dat_rsp_conv_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1437.4]
  wire [7:0] dat_rsp_conv_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1439.4]
  wire [7:0] dat_rsp_conv_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1441.4]
  wire [7:0] dat_rsp_conv_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1443.4]
  wire [7:0] dat_rsp_conv_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1445.4]
  wire [7:0] dat_rsp_conv_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1447.4]
  wire [7:0] dat_rsp_conv_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1449.4]
  wire [7:0] dat_rsp_conv_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1451.4]
  wire [7:0] dat_rsp_conv_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1453.4]
  wire [7:0] dat_rsp_conv_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1455.4]
  wire [7:0] dat_rsp_conv_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1457.4]
  wire [7:0] dat_rsp_conv_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1459.4]
  wire [7:0] dat_rsp_conv_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1461.4]
  wire [7:0] dat_rsp_conv_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1463.4]
  wire [7:0] dat_rsp_conv_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1465.4]
  wire [7:0] dat_rsp_conv_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1467.4]
  wire [7:0] dat_rsp_conv_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1469.4]
  wire [7:0] dat_rsp_conv_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1471.4]
  wire [7:0] dat_rsp_conv_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1473.4]
  wire [7:0] dat_rsp_conv_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1475.4]
  wire [7:0] dat_rsp_conv_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1477.4]
  wire [7:0] dat_rsp_conv_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1479.4]
  wire [7:0] dat_rsp_conv_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1481.4]
  wire [7:0] dat_rsp_conv_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1483.4]
  wire [7:0] dat_rsp_conv_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1485.4]
  wire [7:0] dat_rsp_conv_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1487.4]
  wire [7:0] dat_rsp_conv_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1489.4]
  wire [7:0] dat_rsp_conv_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1491.4]
  wire [7:0] dat_rsp_conv_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1493.4]
  wire [7:0] dat_rsp_conv_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1495.4]
  wire [7:0] dat_rsp_conv_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1497.4]
  wire [7:0] dat_rsp_conv_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1499.4]
  wire [7:0] dat_rsp_conv_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1501.4]
  wire [7:0] dat_rsp_conv_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1503.4]
  wire [7:0] dat_rsp_conv_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1505.4]
  wire [7:0] dat_rsp_conv_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1507.4]
  wire [7:0] dat_rsp_conv_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1509.4]
  wire [7:0] dat_rsp_conv_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1511.4]
  wire [7:0] dat_rsp_conv_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1513.4]
  wire [7:0] dat_rsp_conv_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1515.4]
  wire [7:0] dat_rsp_conv_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1517.4]
  wire [7:0] dat_rsp_conv_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1519.4]
  wire [7:0] dat_rsp_conv_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1521.4]
  wire [7:0] dat_rsp_conv_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1523.4]
  wire [7:0] dat_rsp_conv_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1525.4]
  wire [7:0] dat_rsp_conv_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1527.4]
  wire [7:0] dat_rsp_conv_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1529.4]
  wire [7:0] dat_rsp_conv_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1531.4]
  wire [7:0] dat_rsp_conv_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1533.4]
  wire [7:0] dat_rsp_conv_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1535.4]
  wire [7:0] dat_rsp_conv_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1537.4]
  wire [7:0] dat_rsp_conv_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1539.4]
  wire [7:0] dat_rsp_conv_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1541.4]
  wire [7:0] dat_rsp_conv_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1543.4]
  wire [7:0] dat_rsp_conv_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1545.4]
  wire [7:0] dat_rsp_conv_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1547.4]
  wire [7:0] dat_rsp_conv_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1549.4]
  wire [7:0] dat_rsp_conv_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1551.4]
  reg [255:0] dat_rsp_l0_sft_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 1068:28:@1553.4]
  reg [255:0] _RAND_146;
  reg [127:0] dat_rsp_l0_sft_d2; // @[NV_NVDLA_CSC_dl_for_check.scala 1069:28:@1554.4]
  reg [127:0] _RAND_147;
  reg [127:0] dat_rsp_l0_sft_d3; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:28:@1555.4]
  reg [127:0] _RAND_148;
  reg [127:0] dat_rsp_l1_sft_d2; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:28:@1556.4]
  reg [127:0] _RAND_149;
  reg [127:0] dat_rsp_l1_sft_d3; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:28:@1557.4]
  reg [127:0] _RAND_150;
  reg [127:0] dat_rsp_l2_sft_d3; // @[NV_NVDLA_CSC_dl_for_check.scala 1075:28:@1558.4]
  reg [127:0] _RAND_151;
  wire  _T_1940; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:39:@1559.4]
  wire  _T_1941; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:29:@1560.4]
  wire [1023:0] _T_1943; // @[Cat.scala 30:58:@1561.4]
  wire [1023:0] dat_rsp_l0_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:28:@1562.4]
  wire  _T_1944; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:39:@1563.4]
  wire  _T_1945; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:29:@1564.4]
  wire [1023:0] _T_1947; // @[Cat.scala 30:58:@1565.4]
  wire [1023:0] dat_rsp_l1_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:28:@1566.4]
  wire  _T_1948; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:39:@1567.4]
  wire  _T_1949; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:29:@1568.4]
  wire [1023:0] dat_rsp_l2_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:28:@1570.4]
  wire  _T_1952; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:39:@1571.4]
  wire  _T_1953; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:29:@1572.4]
  wire [1023:0] dat_rsp_l3_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:28:@1574.4]
  wire [10:0] _T_1957; // @[Cat.scala 30:58:@1575.4]
  wire [1023:0] _T_1958; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:41:@1576.4]
  wire [511:0] dat_rsp_l0_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:82:@1577.4]
  wire [10:0] _T_1960; // @[Cat.scala 30:58:@1578.4]
  wire [1023:0] _T_1961; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:41:@1579.4]
  wire [511:0] dat_rsp_l1_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:82:@1580.4]
  wire [10:0] _T_1963; // @[Cat.scala 30:58:@1581.4]
  wire [1023:0] _T_1964; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:41:@1582.4]
  wire [511:0] dat_rsp_l2_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:82:@1583.4]
  wire [10:0] _T_1966; // @[Cat.scala 30:58:@1584.4]
  wire [1023:0] _T_1967; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:41:@1585.4]
  wire [511:0] dat_rsp_l3_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:82:@1586.4]
  wire  _T_1968; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:36:@1587.4]
  wire  _T_1969; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:26:@1588.4]
  wire  _T_1972; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:41:@1589.4]
  wire [127:0] _T_1973; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:81:@1590.4]
  wire [511:0] _T_1979; // @[Cat.scala 30:58:@1596.4]
  wire  _T_1981; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:41:@1597.4]
  wire [255:0] _T_1982; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:81:@1598.4]
  wire [511:0] _T_1984; // @[Cat.scala 30:58:@1600.4]
  wire [511:0] _T_1986; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:25:@1602.4]
  wire [511:0] _T_1987; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:25:@1603.4]
  wire [511:0] dat_rsp_img_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:25:@1604.4]
  wire [7:0] dat_rsp_img_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1606.4]
  wire [7:0] dat_rsp_img_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1608.4]
  wire [7:0] dat_rsp_img_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1610.4]
  wire [7:0] dat_rsp_img_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1612.4]
  wire [7:0] dat_rsp_img_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1614.4]
  wire [7:0] dat_rsp_img_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1616.4]
  wire [7:0] dat_rsp_img_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1618.4]
  wire [7:0] dat_rsp_img_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1620.4]
  wire [7:0] dat_rsp_img_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1622.4]
  wire [7:0] dat_rsp_img_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1624.4]
  wire [7:0] dat_rsp_img_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1626.4]
  wire [7:0] dat_rsp_img_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1628.4]
  wire [7:0] dat_rsp_img_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1630.4]
  wire [7:0] dat_rsp_img_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1632.4]
  wire [7:0] dat_rsp_img_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1634.4]
  wire [7:0] dat_rsp_img_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1636.4]
  wire [7:0] dat_rsp_img_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1638.4]
  wire [7:0] dat_rsp_img_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1640.4]
  wire [7:0] dat_rsp_img_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1642.4]
  wire [7:0] dat_rsp_img_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1644.4]
  wire [7:0] dat_rsp_img_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1646.4]
  wire [7:0] dat_rsp_img_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1648.4]
  wire [7:0] dat_rsp_img_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1650.4]
  wire [7:0] dat_rsp_img_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1652.4]
  wire [7:0] dat_rsp_img_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1654.4]
  wire [7:0] dat_rsp_img_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1656.4]
  wire [7:0] dat_rsp_img_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1658.4]
  wire [7:0] dat_rsp_img_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1660.4]
  wire [7:0] dat_rsp_img_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1662.4]
  wire [7:0] dat_rsp_img_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1664.4]
  wire [7:0] dat_rsp_img_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1666.4]
  wire [7:0] dat_rsp_img_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1668.4]
  wire [7:0] dat_rsp_img_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1670.4]
  wire [7:0] dat_rsp_img_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1672.4]
  wire [7:0] dat_rsp_img_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1674.4]
  wire [7:0] dat_rsp_img_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1676.4]
  wire [7:0] dat_rsp_img_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1678.4]
  wire [7:0] dat_rsp_img_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1680.4]
  wire [7:0] dat_rsp_img_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1682.4]
  wire [7:0] dat_rsp_img_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1684.4]
  wire [7:0] dat_rsp_img_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1686.4]
  wire [7:0] dat_rsp_img_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1688.4]
  wire [7:0] dat_rsp_img_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1690.4]
  wire [7:0] dat_rsp_img_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1692.4]
  wire [7:0] dat_rsp_img_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1694.4]
  wire [7:0] dat_rsp_img_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1696.4]
  wire [7:0] dat_rsp_img_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1698.4]
  wire [7:0] dat_rsp_img_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1700.4]
  wire [7:0] dat_rsp_img_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1702.4]
  wire [7:0] dat_rsp_img_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1704.4]
  wire [7:0] dat_rsp_img_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1706.4]
  wire [7:0] dat_rsp_img_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1708.4]
  wire [7:0] dat_rsp_img_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1710.4]
  wire [7:0] dat_rsp_img_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1712.4]
  wire [7:0] dat_rsp_img_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1714.4]
  wire [7:0] dat_rsp_img_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1716.4]
  wire [7:0] dat_rsp_img_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1718.4]
  wire [7:0] dat_rsp_img_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1720.4]
  wire [7:0] dat_rsp_img_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1722.4]
  wire [7:0] dat_rsp_img_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1724.4]
  wire [7:0] dat_rsp_img_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1726.4]
  wire [7:0] dat_rsp_img_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1728.4]
  wire [7:0] dat_rsp_img_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1730.4]
  wire [7:0] dat_rsp_img_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1732.4]
  wire  _T_2122; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:59:@1734.4]
  wire  dat_rsp_sft_d1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:41:@1735.4]
  wire  _T_2124; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:59:@1736.4]
  wire  dat_rsp_sft_d2_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:41:@1737.4]
  wire  dat_rsp_sft_d3_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:41:@1739.4]
  wire [511:0] _GEN_149; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:24:@1740.4]
  wire [255:0] _GEN_150; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1743.4]
  wire [511:0] _GEN_151; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1743.4]
  wire [511:0] _GEN_154; // @[NV_NVDLA_CSC_dl_for_check.scala 1109:24:@1747.4]
  wire [318:0] _T_2132; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:56:@1753.4]
  wire [63:0] _T_2133; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:73:@1754.4]
  wire [63:0] dat_rsp_ori_mask; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:24:@1755.4]
  wire  _T_2135; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:51:@1756.4]
  wire [63:0] dat_rsp_cur_h_mask_p1; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:32:@1758.4]
  wire  _T_2143; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:51:@1759.4]
  wire [31:0] dat_rsp_cur_h_mask_p2; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:32:@1761.4]
  wire  _T_2151; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:51:@1762.4]
  wire [31:0] dat_rsp_cur_h_mask_p3; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:32:@1764.4]
  wire [31:0] _T_2158; // @[NV_NVDLA_CSC_dl_for_check.scala 1124:57:@1765.4]
  wire [63:0] dat_rsp_cur_h_e2_mask_8b; // @[Cat.scala 30:58:@1767.4]
  wire [15:0] _T_2164; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:57:@1768.4]
  wire [15:0] _T_2165; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:106:@1769.4]
  wire [15:0] _T_2166; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:155:@1770.4]
  wire [63:0] dat_rsp_cur_h_e4_mask_8b; // @[Cat.scala 30:58:@1774.4]
  wire  _T_2175; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:43:@1775.4]
  wire [15:0] _T_2176; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:89:@1776.4]
  wire [63:0] _T_2178; // @[Cat.scala 30:58:@1778.4]
  wire [63:0] _T_2179; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:116:@1779.4]
  wire  _T_2181; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:43:@1780.4]
  wire [31:0] _T_2182; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:89:@1781.4]
  wire [63:0] _T_2183; // @[Cat.scala 30:58:@1782.4]
  wire [63:0] _T_2184; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:116:@1783.4]
  wire [63:0] _T_2185; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:26:@1784.4]
  wire [63:0] dat_rsp_mask_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:26:@1785.4]
  wire  _T_2186; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:35:@1786.4]
  wire [7:0] dat_rsp_data_w_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire [7:0] dat_rsp_data_w_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  wire  dat_rsp_mask_val_int8_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1788.4]
  wire  dat_rsp_mask_val_int8_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1789.4]
  wire  dat_rsp_mask_val_int8_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1790.4]
  wire  dat_rsp_mask_val_int8_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1791.4]
  wire  dat_rsp_mask_val_int8_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1792.4]
  wire  dat_rsp_mask_val_int8_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1793.4]
  wire  dat_rsp_mask_val_int8_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1794.4]
  wire  dat_rsp_mask_val_int8_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1795.4]
  wire  dat_rsp_mask_val_int8_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1796.4]
  wire  dat_rsp_mask_val_int8_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1797.4]
  wire  dat_rsp_mask_val_int8_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1798.4]
  wire  dat_rsp_mask_val_int8_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1799.4]
  wire  dat_rsp_mask_val_int8_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1800.4]
  wire  dat_rsp_mask_val_int8_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1801.4]
  wire  dat_rsp_mask_val_int8_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1802.4]
  wire  dat_rsp_mask_val_int8_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1803.4]
  wire  dat_rsp_mask_val_int8_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1804.4]
  wire  dat_rsp_mask_val_int8_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1805.4]
  wire  dat_rsp_mask_val_int8_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1806.4]
  wire  dat_rsp_mask_val_int8_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1807.4]
  wire  dat_rsp_mask_val_int8_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1808.4]
  wire  dat_rsp_mask_val_int8_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1809.4]
  wire  dat_rsp_mask_val_int8_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1810.4]
  wire  dat_rsp_mask_val_int8_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1811.4]
  wire  dat_rsp_mask_val_int8_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1812.4]
  wire  dat_rsp_mask_val_int8_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1813.4]
  wire  dat_rsp_mask_val_int8_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1814.4]
  wire  dat_rsp_mask_val_int8_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1815.4]
  wire  dat_rsp_mask_val_int8_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1816.4]
  wire  dat_rsp_mask_val_int8_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1817.4]
  wire  dat_rsp_mask_val_int8_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1818.4]
  wire  dat_rsp_mask_val_int8_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1819.4]
  wire  dat_rsp_mask_val_int8_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1820.4]
  wire  dat_rsp_mask_val_int8_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1821.4]
  wire  dat_rsp_mask_val_int8_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1822.4]
  wire  dat_rsp_mask_val_int8_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1823.4]
  wire  dat_rsp_mask_val_int8_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1824.4]
  wire  dat_rsp_mask_val_int8_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1825.4]
  wire  dat_rsp_mask_val_int8_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1826.4]
  wire  dat_rsp_mask_val_int8_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1827.4]
  wire  dat_rsp_mask_val_int8_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1828.4]
  wire  dat_rsp_mask_val_int8_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1829.4]
  wire  dat_rsp_mask_val_int8_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1830.4]
  wire  dat_rsp_mask_val_int8_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1831.4]
  wire  dat_rsp_mask_val_int8_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1832.4]
  wire  dat_rsp_mask_val_int8_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1833.4]
  wire  dat_rsp_mask_val_int8_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1834.4]
  wire  dat_rsp_mask_val_int8_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1835.4]
  wire  dat_rsp_mask_val_int8_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1836.4]
  wire  dat_rsp_mask_val_int8_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1837.4]
  wire  dat_rsp_mask_val_int8_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1838.4]
  wire  dat_rsp_mask_val_int8_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1839.4]
  wire  dat_rsp_mask_val_int8_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1840.4]
  wire  dat_rsp_mask_val_int8_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1841.4]
  wire  dat_rsp_mask_val_int8_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1842.4]
  wire  dat_rsp_mask_val_int8_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1843.4]
  wire  dat_rsp_mask_val_int8_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1844.4]
  wire  dat_rsp_mask_val_int8_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1845.4]
  wire  dat_rsp_mask_val_int8_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1846.4]
  wire  dat_rsp_mask_val_int8_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1847.4]
  wire  dat_rsp_mask_val_int8_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1848.4]
  wire  dat_rsp_mask_val_int8_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1849.4]
  wire  dat_rsp_mask_val_int8_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1850.4]
  wire  dat_rsp_mask_val_int8_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1851.4]
  wire  _T_2515; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1917.4]
  wire  dat_rsp_mask_w_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1918.4]
  wire  _T_2517; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1919.4]
  wire  dat_rsp_mask_w_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1920.4]
  wire  _T_2519; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1921.4]
  wire  dat_rsp_mask_w_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1922.4]
  wire  _T_2521; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1923.4]
  wire  dat_rsp_mask_w_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1924.4]
  wire  _T_2523; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1925.4]
  wire  dat_rsp_mask_w_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1926.4]
  wire  _T_2525; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1927.4]
  wire  dat_rsp_mask_w_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1928.4]
  wire  _T_2527; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1929.4]
  wire  dat_rsp_mask_w_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1930.4]
  wire  _T_2529; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1931.4]
  wire  dat_rsp_mask_w_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1932.4]
  wire  _T_2531; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1933.4]
  wire  dat_rsp_mask_w_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1934.4]
  wire  _T_2533; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1935.4]
  wire  dat_rsp_mask_w_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1936.4]
  wire  _T_2535; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1937.4]
  wire  dat_rsp_mask_w_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1938.4]
  wire  _T_2537; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1939.4]
  wire  dat_rsp_mask_w_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1940.4]
  wire  _T_2539; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1941.4]
  wire  dat_rsp_mask_w_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1942.4]
  wire  _T_2541; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1943.4]
  wire  dat_rsp_mask_w_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1944.4]
  wire  _T_2543; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1945.4]
  wire  dat_rsp_mask_w_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1946.4]
  wire  _T_2545; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1947.4]
  wire  dat_rsp_mask_w_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1948.4]
  wire  _T_2547; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1949.4]
  wire  dat_rsp_mask_w_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1950.4]
  wire  _T_2549; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1951.4]
  wire  dat_rsp_mask_w_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1952.4]
  wire  _T_2551; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1953.4]
  wire  dat_rsp_mask_w_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1954.4]
  wire  _T_2553; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1955.4]
  wire  dat_rsp_mask_w_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1956.4]
  wire  _T_2555; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1957.4]
  wire  dat_rsp_mask_w_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1958.4]
  wire  _T_2557; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1959.4]
  wire  dat_rsp_mask_w_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1960.4]
  wire  _T_2559; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1961.4]
  wire  dat_rsp_mask_w_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1962.4]
  wire  _T_2561; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1963.4]
  wire  dat_rsp_mask_w_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1964.4]
  wire  _T_2563; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1965.4]
  wire  dat_rsp_mask_w_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1966.4]
  wire  _T_2565; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1967.4]
  wire  dat_rsp_mask_w_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1968.4]
  wire  _T_2567; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1969.4]
  wire  dat_rsp_mask_w_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1970.4]
  wire  _T_2569; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1971.4]
  wire  dat_rsp_mask_w_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1972.4]
  wire  _T_2571; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1973.4]
  wire  dat_rsp_mask_w_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1974.4]
  wire  _T_2573; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1975.4]
  wire  dat_rsp_mask_w_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1976.4]
  wire  _T_2575; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1977.4]
  wire  dat_rsp_mask_w_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1978.4]
  wire  _T_2577; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1979.4]
  wire  dat_rsp_mask_w_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1980.4]
  wire  _T_2579; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1981.4]
  wire  dat_rsp_mask_w_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1982.4]
  wire  _T_2581; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1983.4]
  wire  dat_rsp_mask_w_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1984.4]
  wire  _T_2583; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1985.4]
  wire  dat_rsp_mask_w_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1986.4]
  wire  _T_2585; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1987.4]
  wire  dat_rsp_mask_w_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1988.4]
  wire  _T_2587; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1989.4]
  wire  dat_rsp_mask_w_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1990.4]
  wire  _T_2589; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1991.4]
  wire  dat_rsp_mask_w_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1992.4]
  wire  _T_2591; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1993.4]
  wire  dat_rsp_mask_w_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1994.4]
  wire  _T_2593; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1995.4]
  wire  dat_rsp_mask_w_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1996.4]
  wire  _T_2595; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1997.4]
  wire  dat_rsp_mask_w_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1998.4]
  wire  _T_2597; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1999.4]
  wire  dat_rsp_mask_w_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2000.4]
  wire  _T_2599; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2001.4]
  wire  dat_rsp_mask_w_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2002.4]
  wire  _T_2601; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2003.4]
  wire  dat_rsp_mask_w_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2004.4]
  wire  _T_2603; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2005.4]
  wire  dat_rsp_mask_w_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2006.4]
  wire  _T_2605; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2007.4]
  wire  dat_rsp_mask_w_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2008.4]
  wire  _T_2607; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2009.4]
  wire  dat_rsp_mask_w_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2010.4]
  wire  _T_2609; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2011.4]
  wire  dat_rsp_mask_w_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2012.4]
  wire  _T_2611; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2013.4]
  wire  dat_rsp_mask_w_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2014.4]
  wire  _T_2613; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2015.4]
  wire  dat_rsp_mask_w_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2016.4]
  wire  _T_2615; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2017.4]
  wire  dat_rsp_mask_w_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2018.4]
  wire  _T_2617; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2019.4]
  wire  dat_rsp_mask_w_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2020.4]
  wire  _T_2619; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2021.4]
  wire  dat_rsp_mask_w_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2022.4]
  wire  _T_2621; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2023.4]
  wire  dat_rsp_mask_w_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2024.4]
  wire  _T_2623; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2025.4]
  wire  dat_rsp_mask_w_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2026.4]
  wire  _T_2625; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2027.4]
  wire  dat_rsp_mask_w_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2028.4]
  wire  _T_2627; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2029.4]
  wire  dat_rsp_mask_w_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2030.4]
  wire  _T_2629; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2031.4]
  wire  dat_rsp_mask_w_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2032.4]
  wire  _T_2631; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2033.4]
  wire  dat_rsp_mask_w_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2034.4]
  wire  _T_2633; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2035.4]
  wire  dat_rsp_mask_w_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2036.4]
  wire  _T_2635; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2037.4]
  wire  dat_rsp_mask_w_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2038.4]
  wire  _T_2637; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2039.4]
  wire  dat_rsp_mask_w_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2040.4]
  wire  _T_2639; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2041.4]
  wire  dat_rsp_mask_w_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2042.4]
  wire  _T_2641; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2043.4]
  wire  dat_rsp_mask_w_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2044.4]
  reg  dat_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:27:@2110.4]
  reg [31:0] _RAND_152;
  reg [8:0] dat_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1142:27:@2111.4]
  reg [31:0] _RAND_153;
  reg  dat_out_bypass_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_154;
  reg  dat_out_bypass_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_155;
  reg  dat_out_bypass_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_156;
  reg  dat_out_bypass_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_157;
  reg  dat_out_bypass_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_158;
  reg  dat_out_bypass_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_159;
  reg  dat_out_bypass_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_160;
  reg  dat_out_bypass_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_161;
  reg  dat_out_bypass_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_162;
  reg  dat_out_bypass_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_163;
  reg  dat_out_bypass_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_164;
  reg  dat_out_bypass_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_165;
  reg  dat_out_bypass_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_166;
  reg  dat_out_bypass_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_167;
  reg  dat_out_bypass_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_168;
  reg  dat_out_bypass_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_169;
  reg  dat_out_bypass_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_170;
  reg  dat_out_bypass_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_171;
  reg  dat_out_bypass_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_172;
  reg  dat_out_bypass_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_173;
  reg  dat_out_bypass_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_174;
  reg  dat_out_bypass_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_175;
  reg  dat_out_bypass_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_176;
  reg  dat_out_bypass_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_177;
  reg  dat_out_bypass_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_178;
  reg  dat_out_bypass_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_179;
  reg  dat_out_bypass_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_180;
  reg  dat_out_bypass_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_181;
  reg  dat_out_bypass_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_182;
  reg  dat_out_bypass_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_183;
  reg  dat_out_bypass_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_184;
  reg  dat_out_bypass_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_185;
  reg  dat_out_bypass_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_186;
  reg  dat_out_bypass_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_187;
  reg  dat_out_bypass_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_188;
  reg  dat_out_bypass_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_189;
  reg  dat_out_bypass_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_190;
  reg  dat_out_bypass_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_191;
  reg  dat_out_bypass_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_192;
  reg  dat_out_bypass_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_193;
  reg  dat_out_bypass_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_194;
  reg  dat_out_bypass_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_195;
  reg  dat_out_bypass_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_196;
  reg  dat_out_bypass_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_197;
  reg  dat_out_bypass_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_198;
  reg  dat_out_bypass_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_199;
  reg  dat_out_bypass_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_200;
  reg  dat_out_bypass_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_201;
  reg  dat_out_bypass_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_202;
  reg  dat_out_bypass_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_203;
  reg  dat_out_bypass_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_204;
  reg  dat_out_bypass_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_205;
  reg  dat_out_bypass_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_206;
  reg  dat_out_bypass_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_207;
  reg  dat_out_bypass_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_208;
  reg  dat_out_bypass_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_209;
  reg  dat_out_bypass_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_210;
  reg  dat_out_bypass_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_211;
  reg  dat_out_bypass_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_212;
  reg  dat_out_bypass_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_213;
  reg  dat_out_bypass_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_214;
  reg  dat_out_bypass_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_215;
  reg  dat_out_bypass_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_216;
  reg  dat_out_bypass_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1143:34:@2177.4]
  reg [31:0] _RAND_217;
  reg [7:0] dat_out_bypass_data_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_218;
  reg [7:0] dat_out_bypass_data_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_219;
  reg [7:0] dat_out_bypass_data_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_220;
  reg [7:0] dat_out_bypass_data_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_221;
  reg [7:0] dat_out_bypass_data_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_222;
  reg [7:0] dat_out_bypass_data_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_223;
  reg [7:0] dat_out_bypass_data_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_224;
  reg [7:0] dat_out_bypass_data_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_225;
  reg [7:0] dat_out_bypass_data_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_226;
  reg [7:0] dat_out_bypass_data_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_227;
  reg [7:0] dat_out_bypass_data_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_228;
  reg [7:0] dat_out_bypass_data_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_229;
  reg [7:0] dat_out_bypass_data_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_230;
  reg [7:0] dat_out_bypass_data_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_231;
  reg [7:0] dat_out_bypass_data_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_232;
  reg [7:0] dat_out_bypass_data_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_233;
  reg [7:0] dat_out_bypass_data_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_234;
  reg [7:0] dat_out_bypass_data_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_235;
  reg [7:0] dat_out_bypass_data_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_236;
  reg [7:0] dat_out_bypass_data_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_237;
  reg [7:0] dat_out_bypass_data_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_238;
  reg [7:0] dat_out_bypass_data_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_239;
  reg [7:0] dat_out_bypass_data_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_240;
  reg [7:0] dat_out_bypass_data_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_241;
  reg [7:0] dat_out_bypass_data_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_242;
  reg [7:0] dat_out_bypass_data_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_243;
  reg [7:0] dat_out_bypass_data_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_244;
  reg [7:0] dat_out_bypass_data_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_245;
  reg [7:0] dat_out_bypass_data_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_246;
  reg [7:0] dat_out_bypass_data_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_247;
  reg [7:0] dat_out_bypass_data_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_248;
  reg [7:0] dat_out_bypass_data_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_249;
  reg [7:0] dat_out_bypass_data_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_250;
  reg [7:0] dat_out_bypass_data_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_251;
  reg [7:0] dat_out_bypass_data_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_252;
  reg [7:0] dat_out_bypass_data_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_253;
  reg [7:0] dat_out_bypass_data_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_254;
  reg [7:0] dat_out_bypass_data_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_255;
  reg [7:0] dat_out_bypass_data_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_256;
  reg [7:0] dat_out_bypass_data_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_257;
  reg [7:0] dat_out_bypass_data_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_258;
  reg [7:0] dat_out_bypass_data_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_259;
  reg [7:0] dat_out_bypass_data_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_260;
  reg [7:0] dat_out_bypass_data_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_261;
  reg [7:0] dat_out_bypass_data_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_262;
  reg [7:0] dat_out_bypass_data_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_263;
  reg [7:0] dat_out_bypass_data_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_264;
  reg [7:0] dat_out_bypass_data_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_265;
  reg [7:0] dat_out_bypass_data_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_266;
  reg [7:0] dat_out_bypass_data_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_267;
  reg [7:0] dat_out_bypass_data_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_268;
  reg [7:0] dat_out_bypass_data_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_269;
  reg [7:0] dat_out_bypass_data_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_270;
  reg [7:0] dat_out_bypass_data_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_271;
  reg [7:0] dat_out_bypass_data_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_272;
  reg [7:0] dat_out_bypass_data_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_273;
  reg [7:0] dat_out_bypass_data_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_274;
  reg [7:0] dat_out_bypass_data_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_275;
  reg [7:0] dat_out_bypass_data_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_276;
  reg [7:0] dat_out_bypass_data_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_277;
  reg [7:0] dat_out_bypass_data_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_278;
  reg [7:0] dat_out_bypass_data_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_279;
  reg [7:0] dat_out_bypass_data_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_280;
  reg [7:0] dat_out_bypass_data_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1144:30:@2178.4]
  reg [31:0] _RAND_281;
  wire [8:0] _GEN_155; // @[NV_NVDLA_CSC_dl_for_check.scala 1154:21:@2180.4]
  wire  _GEN_156; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_157; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_158; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_159; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_160; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_161; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_162; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_163; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_164; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_165; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_209; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  wire  _T_3247; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2249.4]
  wire  _T_3248; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2253.4]
  wire  _T_3249; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2257.4]
  wire  _T_3250; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2261.4]
  wire  _T_3251; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2265.4]
  wire  _T_3252; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2269.4]
  wire  _T_3253; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2273.4]
  wire  _T_3254; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2277.4]
  wire  _T_3255; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2281.4]
  wire  _T_3256; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2285.4]
  wire  _T_3257; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2289.4]
  wire  _T_3258; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2293.4]
  wire  _T_3259; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2297.4]
  wire  _T_3260; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2301.4]
  wire  _T_3261; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2305.4]
  wire  _T_3262; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2309.4]
  wire  _T_3263; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2313.4]
  wire  _T_3264; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2317.4]
  wire  _T_3265; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2321.4]
  wire  _T_3266; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2325.4]
  wire  _T_3267; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2329.4]
  wire  _T_3268; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2333.4]
  wire  _T_3269; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2337.4]
  wire  _T_3270; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2341.4]
  wire  _T_3271; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2345.4]
  wire  _T_3272; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2349.4]
  wire  _T_3273; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2353.4]
  wire  _T_3274; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2357.4]
  wire  _T_3275; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2361.4]
  wire  _T_3276; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2365.4]
  wire  _T_3277; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2369.4]
  wire  _T_3278; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2373.4]
  wire  _T_3279; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2377.4]
  wire  _T_3280; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2381.4]
  wire  _T_3281; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2385.4]
  wire  _T_3282; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2389.4]
  wire  _T_3283; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2393.4]
  wire  _T_3284; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2397.4]
  wire  _T_3285; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2401.4]
  wire  _T_3286; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2405.4]
  wire  _T_3287; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2409.4]
  wire  _T_3288; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2413.4]
  wire  _T_3289; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2417.4]
  wire  _T_3290; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2421.4]
  wire  _T_3291; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2425.4]
  wire  _T_3292; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2429.4]
  wire  _T_3293; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2433.4]
  wire  _T_3294; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2437.4]
  wire  _T_3295; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2441.4]
  wire  _T_3296; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2445.4]
  wire  _T_3297; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2449.4]
  wire  _T_3298; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2453.4]
  wire  _T_3299; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2457.4]
  wire  _T_3300; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2461.4]
  wire  _T_3301; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2465.4]
  wire  _T_3302; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2469.4]
  wire  _T_3303; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2473.4]
  wire  _T_3304; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2477.4]
  wire  _T_3305; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2481.4]
  wire  _T_3306; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2485.4]
  wire  _T_3307; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2489.4]
  wire  _T_3308; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2493.4]
  wire  _T_3309; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2497.4]
  wire  _T_3310; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2501.4]
  reg  dl_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1169:26:@2505.4]
  reg [31:0] _RAND_282;
  reg  dl_out_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_283;
  reg  dl_out_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_284;
  reg  dl_out_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_285;
  reg  dl_out_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_286;
  reg  dl_out_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_287;
  reg  dl_out_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_288;
  reg  dl_out_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_289;
  reg  dl_out_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_290;
  reg  dl_out_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_291;
  reg  dl_out_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_292;
  reg  dl_out_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_293;
  reg  dl_out_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_294;
  reg  dl_out_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_295;
  reg  dl_out_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_296;
  reg  dl_out_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_297;
  reg  dl_out_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_298;
  reg  dl_out_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_299;
  reg  dl_out_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_300;
  reg  dl_out_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_301;
  reg  dl_out_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_302;
  reg  dl_out_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_303;
  reg  dl_out_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_304;
  reg  dl_out_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_305;
  reg  dl_out_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_306;
  reg  dl_out_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_307;
  reg  dl_out_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_308;
  reg  dl_out_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_309;
  reg  dl_out_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_310;
  reg  dl_out_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_311;
  reg  dl_out_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_312;
  reg  dl_out_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_313;
  reg  dl_out_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_314;
  reg  dl_out_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_315;
  reg  dl_out_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_316;
  reg  dl_out_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_317;
  reg  dl_out_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_318;
  reg  dl_out_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_319;
  reg  dl_out_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_320;
  reg  dl_out_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_321;
  reg  dl_out_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_322;
  reg  dl_out_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_323;
  reg  dl_out_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_324;
  reg  dl_out_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_325;
  reg  dl_out_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_326;
  reg  dl_out_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_327;
  reg  dl_out_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_328;
  reg  dl_out_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_329;
  reg  dl_out_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_330;
  reg  dl_out_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_331;
  reg  dl_out_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_332;
  reg  dl_out_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_333;
  reg  dl_out_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_334;
  reg  dl_out_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_335;
  reg  dl_out_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_336;
  reg  dl_out_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_337;
  reg  dl_out_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_338;
  reg  dl_out_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_339;
  reg  dl_out_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_340;
  reg  dl_out_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_341;
  reg  dl_out_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_342;
  reg  dl_out_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_343;
  reg  dl_out_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_344;
  reg  dl_out_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_345;
  reg  dl_out_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1170:26:@2571.4]
  reg [31:0] _RAND_346;
  reg [8:0] dl_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1171:26:@2572.4]
  reg [31:0] _RAND_347;
  reg [7:0] dl_out_data_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_348;
  reg [7:0] dl_out_data_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_349;
  reg [7:0] dl_out_data_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_350;
  reg [7:0] dl_out_data_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_351;
  reg [7:0] dl_out_data_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_352;
  reg [7:0] dl_out_data_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_353;
  reg [7:0] dl_out_data_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_354;
  reg [7:0] dl_out_data_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_355;
  reg [7:0] dl_out_data_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_356;
  reg [7:0] dl_out_data_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_357;
  reg [7:0] dl_out_data_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_358;
  reg [7:0] dl_out_data_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_359;
  reg [7:0] dl_out_data_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_360;
  reg [7:0] dl_out_data_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_361;
  reg [7:0] dl_out_data_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_362;
  reg [7:0] dl_out_data_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_363;
  reg [7:0] dl_out_data_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_364;
  reg [7:0] dl_out_data_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_365;
  reg [7:0] dl_out_data_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_366;
  reg [7:0] dl_out_data_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_367;
  reg [7:0] dl_out_data_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_368;
  reg [7:0] dl_out_data_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_369;
  reg [7:0] dl_out_data_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_370;
  reg [7:0] dl_out_data_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_371;
  reg [7:0] dl_out_data_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_372;
  reg [7:0] dl_out_data_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_373;
  reg [7:0] dl_out_data_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_374;
  reg [7:0] dl_out_data_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_375;
  reg [7:0] dl_out_data_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_376;
  reg [7:0] dl_out_data_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_377;
  reg [7:0] dl_out_data_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_378;
  reg [7:0] dl_out_data_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_379;
  reg [7:0] dl_out_data_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_380;
  reg [7:0] dl_out_data_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_381;
  reg [7:0] dl_out_data_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_382;
  reg [7:0] dl_out_data_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_383;
  reg [7:0] dl_out_data_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_384;
  reg [7:0] dl_out_data_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_385;
  reg [7:0] dl_out_data_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_386;
  reg [7:0] dl_out_data_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_387;
  reg [7:0] dl_out_data_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_388;
  reg [7:0] dl_out_data_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_389;
  reg [7:0] dl_out_data_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_390;
  reg [7:0] dl_out_data_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_391;
  reg [7:0] dl_out_data_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_392;
  reg [7:0] dl_out_data_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_393;
  reg [7:0] dl_out_data_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_394;
  reg [7:0] dl_out_data_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_395;
  reg [7:0] dl_out_data_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_396;
  reg [7:0] dl_out_data_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_397;
  reg [7:0] dl_out_data_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_398;
  reg [7:0] dl_out_data_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_399;
  reg [7:0] dl_out_data_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_400;
  reg [7:0] dl_out_data_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_401;
  reg [7:0] dl_out_data_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_402;
  reg [7:0] dl_out_data_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_403;
  reg [7:0] dl_out_data_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_404;
  reg [7:0] dl_out_data_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_405;
  reg [7:0] dl_out_data_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_406;
  reg [7:0] dl_out_data_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_407;
  reg [7:0] dl_out_data_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_408;
  reg [7:0] dl_out_data_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_409;
  reg [7:0] dl_out_data_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_410;
  reg [7:0] dl_out_data_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1172:22:@2573.4]
  reg [31:0] _RAND_411;
  wire  _T_3846; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:24:@2574.4]
  wire  dat_out_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  dat_out_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  wire  _T_4112; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:19:@2642.4]
  wire  _GEN_284; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_285; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_286; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_287; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_288; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_289; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_290; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_291; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_292; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_293; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  wire [8:0] _GEN_348; // @[NV_NVDLA_CSC_dl_for_check.scala 1182:19:@2709.4]
  reg  dl_out_pvld_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 1195:29:@2904.4]
  reg [31:0] _RAND_412;
  wire  _T_4115; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:27:@2906.4]
  wire [8:0] sc2mac_dat_pd_w; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:26:@2907.4]
  reg  _T_4119; // @[NV_NVDLA_CSC_dl_for_check.scala 1198:33:@2908.4]
  reg [31:0] _RAND_413;
  reg  _T_4122; // @[NV_NVDLA_CSC_dl_for_check.scala 1199:33:@2911.4]
  reg [31:0] _RAND_414;
  wire  _T_4124; // @[NV_NVDLA_CSC_dl_for_check.scala 1200:85:@2914.4]
  reg [8:0] _T_4126; // @[Reg.scala 19:20:@2915.4]
  reg [31:0] _RAND_415;
  wire [8:0] _GEN_413; // @[Reg.scala 20:19:@2916.4]
  reg [8:0] _T_4130; // @[Reg.scala 19:20:@2921.4]
  reg [31:0] _RAND_416;
  wire [8:0] _GEN_414; // @[Reg.scala 20:19:@2922.4]
  reg  _T_4398_0; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_417;
  reg  _T_4398_1; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_418;
  reg  _T_4398_2; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_419;
  reg  _T_4398_3; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_420;
  reg  _T_4398_4; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_421;
  reg  _T_4398_5; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_422;
  reg  _T_4398_6; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_423;
  reg  _T_4398_7; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_424;
  reg  _T_4398_8; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_425;
  reg  _T_4398_9; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_426;
  reg  _T_4398_10; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_427;
  reg  _T_4398_11; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_428;
  reg  _T_4398_12; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_429;
  reg  _T_4398_13; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_430;
  reg  _T_4398_14; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_431;
  reg  _T_4398_15; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_432;
  reg  _T_4398_16; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_433;
  reg  _T_4398_17; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_434;
  reg  _T_4398_18; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_435;
  reg  _T_4398_19; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_436;
  reg  _T_4398_20; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_437;
  reg  _T_4398_21; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_438;
  reg  _T_4398_22; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_439;
  reg  _T_4398_23; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_440;
  reg  _T_4398_24; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_441;
  reg  _T_4398_25; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_442;
  reg  _T_4398_26; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_443;
  reg  _T_4398_27; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_444;
  reg  _T_4398_28; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_445;
  reg  _T_4398_29; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_446;
  reg  _T_4398_30; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_447;
  reg  _T_4398_31; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_448;
  reg  _T_4398_32; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_449;
  reg  _T_4398_33; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_450;
  reg  _T_4398_34; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_451;
  reg  _T_4398_35; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_452;
  reg  _T_4398_36; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_453;
  reg  _T_4398_37; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_454;
  reg  _T_4398_38; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_455;
  reg  _T_4398_39; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_456;
  reg  _T_4398_40; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_457;
  reg  _T_4398_41; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_458;
  reg  _T_4398_42; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_459;
  reg  _T_4398_43; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_460;
  reg  _T_4398_44; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_461;
  reg  _T_4398_45; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_462;
  reg  _T_4398_46; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_463;
  reg  _T_4398_47; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_464;
  reg  _T_4398_48; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_465;
  reg  _T_4398_49; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_466;
  reg  _T_4398_50; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_467;
  reg  _T_4398_51; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_468;
  reg  _T_4398_52; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_469;
  reg  _T_4398_53; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_470;
  reg  _T_4398_54; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_471;
  reg  _T_4398_55; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_472;
  reg  _T_4398_56; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_473;
  reg  _T_4398_57; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_474;
  reg  _T_4398_58; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_475;
  reg  _T_4398_59; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_476;
  reg  _T_4398_60; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_477;
  reg  _T_4398_61; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_478;
  reg  _T_4398_62; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_479;
  reg  _T_4398_63; // @[Reg.scala 19:20:@2992.4]
  reg [31:0] _RAND_480;
  wire  _GEN_415; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_416; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_417; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_418; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_419; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_420; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_421; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_422; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_423; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_424; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_425; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_426; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_427; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_428; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_429; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_430; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_431; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_432; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_433; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_434; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_435; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_436; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_437; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_438; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_439; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_440; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_441; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_442; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_443; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_444; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_445; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_446; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_447; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_448; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_449; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_450; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_451; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_452; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_453; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_454; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_455; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_456; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_457; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_458; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_459; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_460; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_461; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_462; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_463; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_464; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_465; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_466; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_467; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_468; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_469; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_470; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_471; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_472; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_473; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_474; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_475; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_476; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_477; // @[Reg.scala 20:19:@2993.4]
  wire  _GEN_478; // @[Reg.scala 20:19:@2993.4]
  wire [7:0] _T_4601; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3065.4]
  wire [15:0] _T_4609; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3073.4]
  wire [7:0] _T_4616; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3080.4]
  wire [31:0] _T_4625; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3089.4]
  wire [7:0] _T_4632; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3096.4]
  wire [15:0] _T_4640; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3104.4]
  wire [7:0] _T_4647; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3111.4]
  wire [31:0] _T_4656; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3120.4]
  reg  _T_4925_0; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_481;
  reg  _T_4925_1; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_482;
  reg  _T_4925_2; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_483;
  reg  _T_4925_3; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_484;
  reg  _T_4925_4; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_485;
  reg  _T_4925_5; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_486;
  reg  _T_4925_6; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_487;
  reg  _T_4925_7; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_488;
  reg  _T_4925_8; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_489;
  reg  _T_4925_9; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_490;
  reg  _T_4925_10; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_491;
  reg  _T_4925_11; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_492;
  reg  _T_4925_12; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_493;
  reg  _T_4925_13; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_494;
  reg  _T_4925_14; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_495;
  reg  _T_4925_15; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_496;
  reg  _T_4925_16; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_497;
  reg  _T_4925_17; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_498;
  reg  _T_4925_18; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_499;
  reg  _T_4925_19; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_500;
  reg  _T_4925_20; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_501;
  reg  _T_4925_21; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_502;
  reg  _T_4925_22; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_503;
  reg  _T_4925_23; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_504;
  reg  _T_4925_24; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_505;
  reg  _T_4925_25; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_506;
  reg  _T_4925_26; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_507;
  reg  _T_4925_27; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_508;
  reg  _T_4925_28; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_509;
  reg  _T_4925_29; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_510;
  reg  _T_4925_30; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_511;
  reg  _T_4925_31; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_512;
  reg  _T_4925_32; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_513;
  reg  _T_4925_33; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_514;
  reg  _T_4925_34; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_515;
  reg  _T_4925_35; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_516;
  reg  _T_4925_36; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_517;
  reg  _T_4925_37; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_518;
  reg  _T_4925_38; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_519;
  reg  _T_4925_39; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_520;
  reg  _T_4925_40; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_521;
  reg  _T_4925_41; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_522;
  reg  _T_4925_42; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_523;
  reg  _T_4925_43; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_524;
  reg  _T_4925_44; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_525;
  reg  _T_4925_45; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_526;
  reg  _T_4925_46; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_527;
  reg  _T_4925_47; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_528;
  reg  _T_4925_48; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_529;
  reg  _T_4925_49; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_530;
  reg  _T_4925_50; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_531;
  reg  _T_4925_51; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_532;
  reg  _T_4925_52; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_533;
  reg  _T_4925_53; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_534;
  reg  _T_4925_54; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_535;
  reg  _T_4925_55; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_536;
  reg  _T_4925_56; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_537;
  reg  _T_4925_57; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_538;
  reg  _T_4925_58; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_539;
  reg  _T_4925_59; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_540;
  reg  _T_4925_60; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_541;
  reg  _T_4925_61; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_542;
  reg  _T_4925_62; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_543;
  reg  _T_4925_63; // @[Reg.scala 19:20:@3189.4]
  reg [31:0] _RAND_544;
  wire  _GEN_479; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_480; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_481; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_482; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_483; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_484; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_485; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_486; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_487; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_488; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_489; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_490; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_491; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_492; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_493; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_494; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_495; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_496; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_497; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_498; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_499; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_500; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_501; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_502; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_503; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_504; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_505; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_506; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_507; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_508; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_509; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_510; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_511; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_512; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_513; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_514; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_515; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_516; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_517; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_518; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_519; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_520; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_521; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_522; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_523; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_524; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_525; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_526; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_527; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_528; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_529; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_530; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_531; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_532; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_533; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_534; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_535; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_536; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_537; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_538; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_539; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_540; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_541; // @[Reg.scala 20:19:@3190.4]
  wire  _GEN_542; // @[Reg.scala 20:19:@3190.4]
  wire [7:0] _T_5128; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3262.4]
  wire [15:0] _T_5136; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3270.4]
  wire [7:0] _T_5143; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3277.4]
  wire [31:0] _T_5152; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3286.4]
  wire [7:0] _T_5159; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3293.4]
  wire [15:0] _T_5167; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3301.4]
  wire [7:0] _T_5174; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3308.4]
  wire [31:0] _T_5183; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3317.4]
  reg [7:0] _T_5186; // @[Reg.scala 11:16:@3320.4]
  reg [31:0] _RAND_545;
  reg [7:0] _T_5188; // @[Reg.scala 11:16:@3325.4]
  reg [31:0] _RAND_546;
  reg [7:0] _T_5190; // @[Reg.scala 11:16:@3330.4]
  reg [31:0] _RAND_547;
  reg [7:0] _T_5192; // @[Reg.scala 11:16:@3335.4]
  reg [31:0] _RAND_548;
  reg [7:0] _T_5194; // @[Reg.scala 11:16:@3340.4]
  reg [31:0] _RAND_549;
  reg [7:0] _T_5196; // @[Reg.scala 11:16:@3345.4]
  reg [31:0] _RAND_550;
  reg [7:0] _T_5198; // @[Reg.scala 11:16:@3350.4]
  reg [31:0] _RAND_551;
  reg [7:0] _T_5200; // @[Reg.scala 11:16:@3355.4]
  reg [31:0] _RAND_552;
  reg [7:0] _T_5202; // @[Reg.scala 11:16:@3360.4]
  reg [31:0] _RAND_553;
  reg [7:0] _T_5204; // @[Reg.scala 11:16:@3365.4]
  reg [31:0] _RAND_554;
  reg [7:0] _T_5206; // @[Reg.scala 11:16:@3370.4]
  reg [31:0] _RAND_555;
  reg [7:0] _T_5208; // @[Reg.scala 11:16:@3375.4]
  reg [31:0] _RAND_556;
  reg [7:0] _T_5210; // @[Reg.scala 11:16:@3380.4]
  reg [31:0] _RAND_557;
  reg [7:0] _T_5212; // @[Reg.scala 11:16:@3385.4]
  reg [31:0] _RAND_558;
  reg [7:0] _T_5214; // @[Reg.scala 11:16:@3390.4]
  reg [31:0] _RAND_559;
  reg [7:0] _T_5216; // @[Reg.scala 11:16:@3395.4]
  reg [31:0] _RAND_560;
  reg [7:0] _T_5218; // @[Reg.scala 11:16:@3400.4]
  reg [31:0] _RAND_561;
  reg [7:0] _T_5220; // @[Reg.scala 11:16:@3405.4]
  reg [31:0] _RAND_562;
  reg [7:0] _T_5222; // @[Reg.scala 11:16:@3410.4]
  reg [31:0] _RAND_563;
  reg [7:0] _T_5224; // @[Reg.scala 11:16:@3415.4]
  reg [31:0] _RAND_564;
  reg [7:0] _T_5226; // @[Reg.scala 11:16:@3420.4]
  reg [31:0] _RAND_565;
  reg [7:0] _T_5228; // @[Reg.scala 11:16:@3425.4]
  reg [31:0] _RAND_566;
  reg [7:0] _T_5230; // @[Reg.scala 11:16:@3430.4]
  reg [31:0] _RAND_567;
  reg [7:0] _T_5232; // @[Reg.scala 11:16:@3435.4]
  reg [31:0] _RAND_568;
  reg [7:0] _T_5234; // @[Reg.scala 11:16:@3440.4]
  reg [31:0] _RAND_569;
  reg [7:0] _T_5236; // @[Reg.scala 11:16:@3445.4]
  reg [31:0] _RAND_570;
  reg [7:0] _T_5238; // @[Reg.scala 11:16:@3450.4]
  reg [31:0] _RAND_571;
  reg [7:0] _T_5240; // @[Reg.scala 11:16:@3455.4]
  reg [31:0] _RAND_572;
  reg [7:0] _T_5242; // @[Reg.scala 11:16:@3460.4]
  reg [31:0] _RAND_573;
  reg [7:0] _T_5244; // @[Reg.scala 11:16:@3465.4]
  reg [31:0] _RAND_574;
  reg [7:0] _T_5246; // @[Reg.scala 11:16:@3470.4]
  reg [31:0] _RAND_575;
  reg [7:0] _T_5248; // @[Reg.scala 11:16:@3475.4]
  reg [31:0] _RAND_576;
  reg [7:0] _T_5250; // @[Reg.scala 11:16:@3480.4]
  reg [31:0] _RAND_577;
  reg [7:0] _T_5252; // @[Reg.scala 11:16:@3485.4]
  reg [31:0] _RAND_578;
  reg [7:0] _T_5254; // @[Reg.scala 11:16:@3490.4]
  reg [31:0] _RAND_579;
  reg [7:0] _T_5256; // @[Reg.scala 11:16:@3495.4]
  reg [31:0] _RAND_580;
  reg [7:0] _T_5258; // @[Reg.scala 11:16:@3500.4]
  reg [31:0] _RAND_581;
  reg [7:0] _T_5260; // @[Reg.scala 11:16:@3505.4]
  reg [31:0] _RAND_582;
  reg [7:0] _T_5262; // @[Reg.scala 11:16:@3510.4]
  reg [31:0] _RAND_583;
  reg [7:0] _T_5264; // @[Reg.scala 11:16:@3515.4]
  reg [31:0] _RAND_584;
  reg [7:0] _T_5266; // @[Reg.scala 11:16:@3520.4]
  reg [31:0] _RAND_585;
  reg [7:0] _T_5268; // @[Reg.scala 11:16:@3525.4]
  reg [31:0] _RAND_586;
  reg [7:0] _T_5270; // @[Reg.scala 11:16:@3530.4]
  reg [31:0] _RAND_587;
  reg [7:0] _T_5272; // @[Reg.scala 11:16:@3535.4]
  reg [31:0] _RAND_588;
  reg [7:0] _T_5274; // @[Reg.scala 11:16:@3540.4]
  reg [31:0] _RAND_589;
  reg [7:0] _T_5276; // @[Reg.scala 11:16:@3545.4]
  reg [31:0] _RAND_590;
  reg [7:0] _T_5278; // @[Reg.scala 11:16:@3550.4]
  reg [31:0] _RAND_591;
  reg [7:0] _T_5280; // @[Reg.scala 11:16:@3555.4]
  reg [31:0] _RAND_592;
  reg [7:0] _T_5282; // @[Reg.scala 11:16:@3560.4]
  reg [31:0] _RAND_593;
  reg [7:0] _T_5284; // @[Reg.scala 11:16:@3565.4]
  reg [31:0] _RAND_594;
  reg [7:0] _T_5286; // @[Reg.scala 11:16:@3570.4]
  reg [31:0] _RAND_595;
  reg [7:0] _T_5288; // @[Reg.scala 11:16:@3575.4]
  reg [31:0] _RAND_596;
  reg [7:0] _T_5290; // @[Reg.scala 11:16:@3580.4]
  reg [31:0] _RAND_597;
  reg [7:0] _T_5292; // @[Reg.scala 11:16:@3585.4]
  reg [31:0] _RAND_598;
  reg [7:0] _T_5294; // @[Reg.scala 11:16:@3590.4]
  reg [31:0] _RAND_599;
  reg [7:0] _T_5296; // @[Reg.scala 11:16:@3595.4]
  reg [31:0] _RAND_600;
  reg [7:0] _T_5298; // @[Reg.scala 11:16:@3600.4]
  reg [31:0] _RAND_601;
  reg [7:0] _T_5300; // @[Reg.scala 11:16:@3605.4]
  reg [31:0] _RAND_602;
  reg [7:0] _T_5302; // @[Reg.scala 11:16:@3610.4]
  reg [31:0] _RAND_603;
  reg [7:0] _T_5304; // @[Reg.scala 11:16:@3615.4]
  reg [31:0] _RAND_604;
  reg [7:0] _T_5306; // @[Reg.scala 11:16:@3620.4]
  reg [31:0] _RAND_605;
  reg [7:0] _T_5308; // @[Reg.scala 11:16:@3625.4]
  reg [31:0] _RAND_606;
  reg [7:0] _T_5310; // @[Reg.scala 11:16:@3630.4]
  reg [31:0] _RAND_607;
  reg [7:0] _T_5312; // @[Reg.scala 11:16:@3635.4]
  reg [31:0] _RAND_608;
  reg [7:0] _T_5314; // @[Reg.scala 11:16:@3640.4]
  reg [31:0] _RAND_609;
  reg [7:0] _T_5316; // @[Reg.scala 11:16:@3645.4]
  reg [31:0] _RAND_610;
  reg [7:0] _T_5318; // @[Reg.scala 11:16:@3650.4]
  reg [31:0] _RAND_611;
  reg [7:0] _T_5320; // @[Reg.scala 11:16:@3655.4]
  reg [31:0] _RAND_612;
  reg [7:0] _T_5322; // @[Reg.scala 11:16:@3660.4]
  reg [31:0] _RAND_613;
  reg [7:0] _T_5324; // @[Reg.scala 11:16:@3665.4]
  reg [31:0] _RAND_614;
  reg [7:0] _T_5326; // @[Reg.scala 11:16:@3670.4]
  reg [31:0] _RAND_615;
  reg [7:0] _T_5328; // @[Reg.scala 11:16:@3675.4]
  reg [31:0] _RAND_616;
  reg [7:0] _T_5330; // @[Reg.scala 11:16:@3680.4]
  reg [31:0] _RAND_617;
  reg [7:0] _T_5332; // @[Reg.scala 11:16:@3685.4]
  reg [31:0] _RAND_618;
  reg [7:0] _T_5334; // @[Reg.scala 11:16:@3690.4]
  reg [31:0] _RAND_619;
  reg [7:0] _T_5336; // @[Reg.scala 11:16:@3695.4]
  reg [31:0] _RAND_620;
  reg [7:0] _T_5338; // @[Reg.scala 11:16:@3700.4]
  reg [31:0] _RAND_621;
  reg [7:0] _T_5340; // @[Reg.scala 11:16:@3705.4]
  reg [31:0] _RAND_622;
  reg [7:0] _T_5342; // @[Reg.scala 11:16:@3710.4]
  reg [31:0] _RAND_623;
  reg [7:0] _T_5344; // @[Reg.scala 11:16:@3715.4]
  reg [31:0] _RAND_624;
  reg [7:0] _T_5346; // @[Reg.scala 11:16:@3720.4]
  reg [31:0] _RAND_625;
  reg [7:0] _T_5348; // @[Reg.scala 11:16:@3725.4]
  reg [31:0] _RAND_626;
  reg [7:0] _T_5350; // @[Reg.scala 11:16:@3730.4]
  reg [31:0] _RAND_627;
  reg [7:0] _T_5352; // @[Reg.scala 11:16:@3735.4]
  reg [31:0] _RAND_628;
  reg [7:0] _T_5354; // @[Reg.scala 11:16:@3740.4]
  reg [31:0] _RAND_629;
  reg [7:0] _T_5356; // @[Reg.scala 11:16:@3745.4]
  reg [31:0] _RAND_630;
  reg [7:0] _T_5358; // @[Reg.scala 11:16:@3750.4]
  reg [31:0] _RAND_631;
  reg [7:0] _T_5360; // @[Reg.scala 11:16:@3755.4]
  reg [31:0] _RAND_632;
  reg [7:0] _T_5362; // @[Reg.scala 11:16:@3760.4]
  reg [31:0] _RAND_633;
  reg [7:0] _T_5364; // @[Reg.scala 11:16:@3765.4]
  reg [31:0] _RAND_634;
  reg [7:0] _T_5366; // @[Reg.scala 11:16:@3770.4]
  reg [31:0] _RAND_635;
  reg [7:0] _T_5368; // @[Reg.scala 11:16:@3775.4]
  reg [31:0] _RAND_636;
  reg [7:0] _T_5370; // @[Reg.scala 11:16:@3780.4]
  reg [31:0] _RAND_637;
  reg [7:0] _T_5372; // @[Reg.scala 11:16:@3785.4]
  reg [31:0] _RAND_638;
  reg [7:0] _T_5374; // @[Reg.scala 11:16:@3790.4]
  reg [31:0] _RAND_639;
  reg [7:0] _T_5376; // @[Reg.scala 11:16:@3795.4]
  reg [31:0] _RAND_640;
  reg [7:0] _T_5378; // @[Reg.scala 11:16:@3800.4]
  reg [31:0] _RAND_641;
  reg [7:0] _T_5380; // @[Reg.scala 11:16:@3805.4]
  reg [31:0] _RAND_642;
  reg [7:0] _T_5382; // @[Reg.scala 11:16:@3810.4]
  reg [31:0] _RAND_643;
  reg [7:0] _T_5384; // @[Reg.scala 11:16:@3815.4]
  reg [31:0] _RAND_644;
  reg [7:0] _T_5386; // @[Reg.scala 11:16:@3820.4]
  reg [31:0] _RAND_645;
  reg [7:0] _T_5388; // @[Reg.scala 11:16:@3825.4]
  reg [31:0] _RAND_646;
  reg [7:0] _T_5390; // @[Reg.scala 11:16:@3830.4]
  reg [31:0] _RAND_647;
  reg [7:0] _T_5392; // @[Reg.scala 11:16:@3835.4]
  reg [31:0] _RAND_648;
  reg [7:0] _T_5394; // @[Reg.scala 11:16:@3840.4]
  reg [31:0] _RAND_649;
  reg [7:0] _T_5396; // @[Reg.scala 11:16:@3845.4]
  reg [31:0] _RAND_650;
  reg [7:0] _T_5398; // @[Reg.scala 11:16:@3850.4]
  reg [31:0] _RAND_651;
  reg [7:0] _T_5400; // @[Reg.scala 11:16:@3855.4]
  reg [31:0] _RAND_652;
  reg [7:0] _T_5402; // @[Reg.scala 11:16:@3860.4]
  reg [31:0] _RAND_653;
  reg [7:0] _T_5404; // @[Reg.scala 11:16:@3865.4]
  reg [31:0] _RAND_654;
  reg [7:0] _T_5406; // @[Reg.scala 11:16:@3870.4]
  reg [31:0] _RAND_655;
  reg [7:0] _T_5408; // @[Reg.scala 11:16:@3875.4]
  reg [31:0] _RAND_656;
  reg [7:0] _T_5410; // @[Reg.scala 11:16:@3880.4]
  reg [31:0] _RAND_657;
  reg [7:0] _T_5412; // @[Reg.scala 11:16:@3885.4]
  reg [31:0] _RAND_658;
  reg [7:0] _T_5414; // @[Reg.scala 11:16:@3890.4]
  reg [31:0] _RAND_659;
  reg [7:0] _T_5416; // @[Reg.scala 11:16:@3895.4]
  reg [31:0] _RAND_660;
  reg [7:0] _T_5418; // @[Reg.scala 11:16:@3900.4]
  reg [31:0] _RAND_661;
  reg [7:0] _T_5420; // @[Reg.scala 11:16:@3905.4]
  reg [31:0] _RAND_662;
  reg [7:0] _T_5422; // @[Reg.scala 11:16:@3910.4]
  reg [31:0] _RAND_663;
  reg [7:0] _T_5424; // @[Reg.scala 11:16:@3915.4]
  reg [31:0] _RAND_664;
  reg [7:0] _T_5426; // @[Reg.scala 11:16:@3920.4]
  reg [31:0] _RAND_665;
  reg [7:0] _T_5428; // @[Reg.scala 11:16:@3925.4]
  reg [31:0] _RAND_666;
  reg [7:0] _T_5430; // @[Reg.scala 11:16:@3930.4]
  reg [31:0] _RAND_667;
  reg [7:0] _T_5432; // @[Reg.scala 11:16:@3935.4]
  reg [31:0] _RAND_668;
  reg [7:0] _T_5434; // @[Reg.scala 11:16:@3940.4]
  reg [31:0] _RAND_669;
  reg [7:0] _T_5436; // @[Reg.scala 11:16:@3945.4]
  reg [31:0] _RAND_670;
  reg [7:0] _T_5438; // @[Reg.scala 11:16:@3950.4]
  reg [31:0] _RAND_671;
  reg [7:0] _T_5440; // @[Reg.scala 11:16:@3955.4]
  reg [31:0] _RAND_672;
  assign _T_337 = nvdla_core_rstn == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 95:38:@8.4]
  assign is_sg_idle = sc_state == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 99:31:@9.4]
  assign is_sg_done = sc_state == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 101:31:@11.4]
  assign layer_st = reg2dp_op_en & is_sg_idle; // @[NV_NVDLA_CSC_dl_for_check.scala 108:32:@14.4]
  assign is_conv = reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 110:35:@16.4]
  assign is_img = is_conv & reg2dp_datain_format; // @[NV_NVDLA_CSC_dl_for_check.scala 111:22:@17.4]
  assign _T_346 = 7'h9 << reg2dp_y_extension; // @[NV_NVDLA_CSC_dl_for_check.scala 118:53:@18.4]
  assign _T_348 = is_img ? _T_346 : 7'h8; // @[NV_NVDLA_CSC_dl_for_check.scala 118:24:@19.4]
  assign sub_h_total_w = _T_348[5:3]; // @[NV_NVDLA_CSC_dl_for_check.scala 118:100:@20.4]
  assign sub_h_cmp_w = is_img ? sub_h_total_w : 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 119:22:@21.4]
  assign _T_351 = sub_h_cmp_w - 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@22.4]
  assign dataout_w_init = $unsigned(_T_351); // @[NV_NVDLA_CSC_dl_for_check.scala 120:34:@23.4]
  assign conv_x_stride_w = reg2dp_conv_x_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 121:51:@24.4]
  assign _T_353 = reg2dp_datain_channel_ext[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 122:62:@25.4]
  assign _T_356 = {conv_x_stride_w,2'h0}; // @[Cat.scala 30:58:@26.4]
  assign _T_359 = {conv_x_stride_w,1'h0}; // @[Cat.scala 30:58:@27.4]
  assign _GEN_671 = {{1'd0}, conv_x_stride_w}; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  assign _T_360 = _T_359 + _GEN_671; // @[NV_NVDLA_CSC_dl_for_check.scala 124:74:@28.4]
  assign _T_361 = 2'h2 == _T_353; // @[Mux.scala 46:19:@29.4]
  assign _T_362 = _T_361 ? _T_360 : {{2'd0}, conv_x_stride_w}; // @[Mux.scala 46:16:@30.4]
  assign _T_363 = 2'h3 == _T_353; // @[Mux.scala 46:19:@31.4]
  assign pixel_x_stride_w = _T_363 ? _T_356 : _T_362; // @[Mux.scala 46:16:@32.4]
  assign _T_365 = reg2dp_weight_channel_ext >= 13'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 126:88:@33.4]
  assign _T_371 = reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 126:172:@35.4]
  assign _T_372 = _T_365 ? 6'h3f : _T_371; // @[NV_NVDLA_CSC_dl_for_check.scala 126:58:@36.4]
  assign _T_375 = {pixel_x_stride_w,1'h0}; // @[Cat.scala 30:58:@37.4]
  assign _GEN_672 = {{1'd0}, pixel_x_stride_w}; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  assign _T_376 = _T_375 + _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@38.4]
  assign _T_377 = _T_375 + _GEN_672; // @[NV_NVDLA_CSC_dl_for_check.scala 127:81:@39.4]
  assign _GEN_673 = {{1'd0}, _T_371}; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  assign _T_379 = _T_377 + _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@41.4]
  assign _T_380 = _T_377 + _GEN_673; // @[NV_NVDLA_CSC_dl_for_check.scala 127:100:@42.4]
  assign _T_383 = pixel_x_stride_w + _T_371; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@44.4]
  assign _T_384 = pixel_x_stride_w + _T_371; // @[NV_NVDLA_CSC_dl_for_check.scala 128:58:@45.4]
  assign _T_385 = 2'h1 == reg2dp_y_extension; // @[Mux.scala 46:19:@46.4]
  assign _T_386 = _T_385 ? _T_384 : _T_372; // @[Mux.scala 46:16:@47.4]
  assign _T_387 = 2'h2 == reg2dp_y_extension; // @[Mux.scala 46:19:@48.4]
  assign pixel_x_init_w = _T_387 ? _T_380 : {{1'd0}, _T_386}; // @[Mux.scala 46:16:@49.4]
  assign pixel_x_init_offset_w = _T_371 + 6'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 129:80:@51.4]
  assign _T_392 = {pixel_x_stride_w,2'h0}; // @[Cat.scala 30:58:@52.4]
  assign _T_397 = _T_385 ? _T_375 : {{1'd0}, pixel_x_stride_w}; // @[Mux.scala 46:16:@55.4]
  assign pixel_x_add_w = _T_387 ? _T_392 : {{1'd0}, _T_397}; // @[Mux.scala 46:16:@57.4]
  assign pixel_ch_stride_w = {pixel_x_stride_w,6'h0}; // @[Cat.scala 30:58:@58.4]
  assign conv_y_stride_w = reg2dp_conv_y_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 139:52:@59.4]
  assign _T_403 = reg2dp_x_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 140:60:@60.4]
  assign x_dilate_w = is_img ? 6'h1 : _T_403; // @[NV_NVDLA_CSC_dl_for_check.scala 140:21:@61.4]
  assign _T_406 = reg2dp_y_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 141:60:@62.4]
  assign y_dilate_w = is_img ? 6'h1 : _T_406; // @[NV_NVDLA_CSC_dl_for_check.scala 141:21:@63.4]
  assign entries_single_w = reg2dp_entries + 14'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 157:43:@87.4]
  assign _T_477 = entries_single_w * 15'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 158:41:@89.4]
  assign entries_batch_w = _T_477[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 158:56:@90.4]
  assign h_offset_slice_w = 6'h1 * y_dilate_w; // @[NV_NVDLA_CSC_dl_for_check.scala 160:37:@91.4]
  assign _GEN_674 = {{9'd0}, data_batch}; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  assign _T_478 = entries * _GEN_674; // @[NV_NVDLA_CSC_dl_for_check.scala 161:34:@92.4]
  assign h_bias_0_stride_w = _T_478[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 161:47:@93.4]
  assign _GEN_675 = {{1'd0}, h_offset_slice}; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  assign _T_479 = entries * _GEN_675; // @[NV_NVDLA_CSC_dl_for_check.scala 162:34:@94.4]
  assign h_bias_1_stride_w = _T_479[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 162:51:@95.4]
  assign rls_slices_w = reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 163:41:@96.4]
  assign _T_482 = reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 164:77:@97.4]
  assign _GEN_676 = {{1'd0}, reg2dp_rls_slices}; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@98.4]
  assign _T_483 = reg2dp_datain_height_ext - _GEN_676; // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@98.4]
  assign _T_484 = $unsigned(_T_483); // @[NV_NVDLA_CSC_dl_for_check.scala 164:113:@99.4]
  assign slice_left_w = reg2dp_skip_data_rls ? _T_482 : _T_484; // @[NV_NVDLA_CSC_dl_for_check.scala 164:23:@100.4]
  assign slices_oprand = layer_st_d1 ? rls_slices : slice_left; // @[NV_NVDLA_CSC_dl_for_check.scala 165:24:@101.4]
  assign _GEN_677 = {{1'd0}, slices_oprand}; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@102.4]
  assign _T_485 = entries_batch * _GEN_677; // @[NV_NVDLA_CSC_dl_for_check.scala 166:38:@102.4]
  assign slice_entries_w = _T_485[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 166:54:@103.4]
  assign _T_670 = is_img ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@174.6]
  assign _T_672 = reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@176.6]
  assign _T_673 = reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 215:38:@177.6]
  assign _T_675 = reg2dp_datain_width_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 216:48:@179.6]
  assign _T_681 = reg2dp_weight_channel_ext[12:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 219:93:@184.6]
  assign _T_682 = {4'h0,_T_681}; // @[Cat.scala 30:58:@185.6]
  assign _T_686 = {1'h0,reg2dp_entries}; // @[Cat.scala 30:58:@218.6]
  assign _GEN_1 = layer_st ? _T_670 : is_img_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_2 = layer_st ? _T_673 : data_bank; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_3 = layer_st ? _T_675 : datain_width; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_4 = layer_st ? reg2dp_datain_width_ext : datain_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_5 = layer_st ? reg2dp_datain_height_ext : datain_height_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_6 = layer_st ? _T_682 : datain_channel_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_7 = layer_st ? sub_h_total_w : sub_h_total_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_8 = layer_st ? sub_h_total_w : sub_h_total_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_10 = layer_st ? sub_h_total_w : sub_h_total_g3; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_11 = layer_st ? sub_h_total_w : sub_h_total_g4; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_12 = layer_st ? sub_h_total_w : sub_h_total_g5; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_13 = layer_st ? sub_h_total_w : sub_h_total_g6; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_15 = layer_st ? sub_h_total_w : sub_h_total_g8; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_16 = layer_st ? sub_h_total_w : sub_h_total_g9; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_18 = layer_st ? sub_h_total_w : sub_h_total_g11; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_19 = layer_st ? sub_h_cmp_w : sub_h_cmp_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_20 = layer_st ? sub_h_cmp_w : sub_h_cmp_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_21 = layer_st ? conv_x_stride_w : conv_x_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_22 = layer_st ? conv_y_stride_w : conv_y_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_24 = layer_st ? 6'h1 : data_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_25 = layer_st ? 5'h0 : batch_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_26 = layer_st ? pixel_x_init_w : pixel_x_init; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_27 = layer_st ? pixel_x_init_offset_w : pixel_x_init_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_28 = layer_st ? pixel_x_add_w : pixel_x_add; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_29 = layer_st ? {{1'd0}, pixel_x_stride_w} : pixel_x_byte_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_30 = layer_st ? pixel_ch_stride_w : pixel_ch_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_31 = layer_st ? x_dilate_w : x_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_32 = layer_st ? y_dilate_w : y_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_33 = layer_st ? reg2dp_pad_value : pad_value; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_34 = layer_st ? entries_single_w : entries; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_35 = layer_st ? entries_batch_w : entries_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_36 = layer_st ? _T_686 : entries_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_37 = layer_st ? {{2'd0}, h_offset_slice_w} : h_offset_slice; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_38 = layer_st ? {{1'd0}, rls_slices_w} : rls_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_39 = layer_st ? slice_left_w : slice_left; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_40 = layer_st ? reg2dp_dataout_width : dataout_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 212:15:@170.4]
  assign _GEN_43 = layer_st_d1 ? h_bias_0_stride_w : h_bias_0_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  assign _GEN_44 = layer_st_d1 ? h_bias_1_stride_w : h_bias_1_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  assign _GEN_45 = layer_st_d1 ? entries : h_bias_2_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  assign _GEN_46 = layer_st_d1 ? entries : h_bias_3_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  assign _GEN_47 = layer_st_d1 ? slice_entries_w : rls_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 257:18:@231.4]
  assign _GEN_48 = is_sg_done ? slice_left : last_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@238.4]
  assign _GEN_49 = is_sg_done ? slice_entries_w : last_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 264:17:@238.4]
  assign _T_763 = last_slices != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 328:37:@313.4]
  assign _T_764 = sg2dl_reuse_rls & _T_763; // @[NV_NVDLA_CSC_dl_for_check.scala 328:23:@314.4]
  assign _T_1627 = sub_h_total_g3[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 918:32:@1216.4]
  assign _T_1628 = _T_1627 & dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 918:36:@1217.4]
  assign _T_1629 = sub_h_total_g3[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 919:35:@1218.4]
  assign _T_1630 = _T_1629 & dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 919:39:@1219.4]
  assign _T_1631 = _T_1628 | _T_1630; // @[NV_NVDLA_CSC_dl_for_check.scala 918:57:@1220.4]
  assign _T_1632 = sub_h_total_g3[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 920:35:@1221.4]
  assign _T_1633 = _T_1632 & dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 920:39:@1222.4]
  assign dat_rsp_pvld = _T_1631 | _T_1633; // @[NV_NVDLA_CSC_dl_for_check.scala 919:60:@1223.4]
  assign _T_1635 = sub_h_total_g4[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 927:42:@1225.4]
  assign _T_1639 = _T_1635 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1227.4]
  assign _T_1640 = _T_1639 & _T_1617; // @[NV_NVDLA_CSC_dl_for_check.scala 927:47:@1228.4]
  assign _T_1641 = sub_h_total_g4[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 928:42:@1229.4]
  assign _T_1645 = _T_1641 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1231.4]
  assign _T_1646 = _T_1645 & _T_1611; // @[NV_NVDLA_CSC_dl_for_check.scala 928:47:@1232.4]
  assign _T_1647 = _T_1640 | _T_1646; // @[NV_NVDLA_CSC_dl_for_check.scala 927:66:@1233.4]
  assign _T_1648 = sub_h_total_g4[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 929:42:@1234.4]
  assign _T_1652 = _T_1648 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1236.4]
  assign _T_1653 = _T_1652 & _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 929:47:@1237.4]
  assign dat_rsp_pd = _T_1647 | _T_1653; // @[NV_NVDLA_CSC_dl_for_check.scala 928:66:@1238.4]
  assign dat_rsp_rls = dat_rsp_pd[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 953:26:@1257.4]
  assign sub_rls = dat_rsp_pvld & dat_rsp_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 325:29:@312.4]
  assign _T_766 = rls_slices != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 328:66:@315.4]
  assign _T_767 = sub_rls & _T_766; // @[NV_NVDLA_CSC_dl_for_check.scala 328:53:@316.4]
  assign dat_rls = _T_764 | _T_767; // @[NV_NVDLA_CSC_dl_for_check.scala 328:42:@317.4]
  assign sc2cdma_dat_slices_w = sub_rls ? rls_slices : last_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 329:28:@319.4]
  assign sc2cdma_dat_entries_w = sub_rls ? rls_entries : last_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 330:29:@321.4]
  assign dat_entry_avl_sub = dat_rls ? sc2cdma_dat_entries_w : 15'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 297:28:@261.4]
  assign _T_720 = dat_entry_st + dat_entry_avl_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@268.4]
  assign dat_entry_st_inc = dat_entry_st + dat_entry_avl_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 302:37:@269.4]
  assign _T_726 = {data_bank,9'h0}; // @[Cat.scala 30:58:@271.4]
  assign _GEN_678 = {{1'd0}, _T_726}; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@272.4]
  assign _T_727 = dat_entry_st_inc - _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@272.4]
  assign _T_728 = $unsigned(_T_727); // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@273.4]
  assign dat_entry_st_inc_wrap = _T_728[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 303:46:@274.4]
  assign is_dat_entry_st_wrap = dat_entry_st_inc >= _GEN_678; // @[NV_NVDLA_CSC_dl_for_check.scala 304:45:@277.4]
  assign _T_736 = is_dat_entry_st_wrap ? dat_entry_st_inc_wrap : dat_entry_st_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 305:83:@278.4]
  assign dat_entry_st_w = sc2cdma_dat_pending_req ? 15'h0 : _T_736; // @[NV_NVDLA_CSC_dl_for_check.scala 305:25:@279.4]
  assign _T_758 = dat_rls | sc2cdma_dat_pending_req; // @[NV_NVDLA_CSC_dl_for_check.scala 316:13:@302.4]
  assign _GEN_52 = _T_758 ? dat_entry_st_w : dat_entry_st; // @[NV_NVDLA_CSC_dl_for_check.scala 316:25:@303.4]
  assign _GEN_54 = dat_rls ? sc2cdma_dat_slices_w : _T_776; // @[Reg.scala 20:19:@327.4]
  assign _GEN_55 = dat_rls ? sc2cdma_dat_entries_w : _T_779; // @[Reg.scala 20:19:@332.4]
  assign _T_828 = {{30'd0}, dl_in_pvld}; // @[NV_NVDLA_CSC_dl_for_check.scala 365:19:@375.4 NV_NVDLA_CSC_dl_for_check.scala 369:12:@381.4]
  assign _GEN_61 = dl_in_pvld ? _T_828 : _T_831; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@383.4]
  assign _GEN_62 = _T_817 ? _T_831 : _T_834; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@387.4]
  assign _GEN_63 = _T_820 ? _T_834 : _T_837; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@391.4]
  assign _GEN_64 = _T_823 ? _T_837 : _T_840; // @[NV_NVDLA_CSC_dl_for_check.scala 373:23:@395.4]
  assign _T_841 = sub_h_total_g0[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 378:30:@398.4]
  assign _T_842 = _T_841 & _T_817; // @[NV_NVDLA_CSC_dl_for_check.scala 378:34:@399.4]
  assign _T_843 = sub_h_total_g0[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 379:30:@400.4]
  assign _T_844 = _T_843 & _T_823; // @[NV_NVDLA_CSC_dl_for_check.scala 379:34:@401.4]
  assign _T_845 = _T_842 | _T_844; // @[NV_NVDLA_CSC_dl_for_check.scala 378:50:@402.4]
  assign _T_846 = sub_h_total_g0[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 380:30:@403.4]
  assign _T_847 = _T_846 & _T_826; // @[NV_NVDLA_CSC_dl_for_check.scala 380:34:@404.4]
  assign dl_pvld = _T_845 | _T_847; // @[NV_NVDLA_CSC_dl_for_check.scala 379:50:@405.4]
  assign _T_848 = sub_h_total_g1[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 382:37:@406.4]
  assign _T_852 = _T_848 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@408.4]
  assign _T_853 = _T_852 & _T_831; // @[NV_NVDLA_CSC_dl_for_check.scala 382:42:@409.4]
  assign _T_854 = sub_h_total_g1[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 383:37:@410.4]
  assign _T_858 = _T_854 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@412.4]
  assign _T_859 = _T_858 & _T_837; // @[NV_NVDLA_CSC_dl_for_check.scala 383:42:@413.4]
  assign _T_860 = _T_853 | _T_859; // @[NV_NVDLA_CSC_dl_for_check.scala 382:56:@414.4]
  assign _T_861 = sub_h_total_g1[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 384:37:@415.4]
  assign _T_865 = _T_861 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@417.4]
  assign _T_866 = _T_865 & _T_840; // @[NV_NVDLA_CSC_dl_for_check.scala 384:42:@418.4]
  assign dl_pd = _T_860 | _T_866; // @[NV_NVDLA_CSC_dl_for_check.scala 383:56:@419.4]
  assign dl_w_offset = dl_pd[4:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 387:24:@420.4]
  assign dl_h_offset = dl_pd[9:5]; // @[NV_NVDLA_CSC_dl_for_check.scala 388:24:@421.4]
  assign dl_channel_size = dl_pd[16:10]; // @[NV_NVDLA_CSC_dl_for_check.scala 389:28:@422.4]
  assign dl_stripe_length = dl_pd[23:17]; // @[NV_NVDLA_CSC_dl_for_check.scala 390:29:@423.4]
  assign dl_cur_sub_h = dl_pd[25:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 391:25:@424.4]
  assign dl_block_end = dl_pd[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 392:25:@425.4]
  assign dl_channel_end = dl_pd[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 393:27:@426.4]
  assign dl_group_end = dl_pd[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 394:25:@427.4]
  assign dl_layer_end = dl_pd[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 395:25:@428.4]
  assign dl_dat_release = dl_pd[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 396:27:@429.4]
  assign _T_874 = batch_cnt + 6'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 405:24:@433.4]
  assign _GEN_682 = {{1'd0}, batch_cmp}; // @[NV_NVDLA_CSC_dl_for_check.scala 407:27:@438.4]
  assign is_batch_end = batch_cnt == _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 407:27:@438.4]
  assign _T_875 = is_batch_end ? 7'h0 : _T_874; // @[NV_NVDLA_CSC_dl_for_check.scala 404:17:@434.4]
  assign _T_876 = layer_st ? 7'h0 : _T_875; // @[NV_NVDLA_CSC_dl_for_check.scala 403:17:@435.4]
  assign _T_877 = _T_876[5:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 405:32:@436.4]
  assign sub_h_cnt_inc = sub_h_cnt + 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 413:31:@442.4]
  assign is_sub_h_end = sub_h_cnt_inc == sub_h_cmp_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 414:32:@443.4]
  assign _T_885 = reg2dp_y_extension != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 415:61:@445.4]
  assign _T_921 = stripe_cnt != 7'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 448:37:@482.4]
  assign _T_922 = ~ _T_921; // @[NV_NVDLA_CSC_dl_for_check.scala 448:24:@483.4]
  assign _T_924 = sub_h_cnt != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 448:56:@484.4]
  assign _T_925 = ~ _T_924; // @[NV_NVDLA_CSC_dl_for_check.scala 448:44:@485.4]
  assign _T_926 = _T_922 & _T_925; // @[NV_NVDLA_CSC_dl_for_check.scala 448:42:@486.4]
  assign _T_928 = batch_cnt != 6'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 448:75:@487.4]
  assign _T_929 = ~ _T_928; // @[NV_NVDLA_CSC_dl_for_check.scala 448:63:@488.4]
  assign _T_930 = _T_926 & _T_929; // @[NV_NVDLA_CSC_dl_for_check.scala 448:61:@489.4]
  assign _T_932 = _T_930 ? 1'h0 : dat_exec_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 448:22:@490.4]
  assign dat_exec_valid = dl_pvld ? 1'h1 : _T_932; // @[NV_NVDLA_CSC_dl_for_check.scala 447:22:@491.4]
  assign _T_886 = _T_885 & dat_exec_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 415:66:@446.4]
  assign sub_h_cnt_reg_en = layer_st | _T_886; // @[NV_NVDLA_CSC_dl_for_check.scala 415:33:@447.4]
  assign _T_887 = layer_st | is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 417:31:@449.6]
  assign _T_889 = _T_887 ? 3'h0 : sub_h_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 417:21:@450.6]
  assign _GEN_65 = sub_h_cnt_reg_en ? _T_889 : {{1'd0}, sub_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 416:23:@448.4]
  assign stripe_cnt_inc = stripe_cnt + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 425:33:@456.4]
  assign _GEN_683 = {{1'd0}, dl_stripe_length}; // @[NV_NVDLA_CSC_dl_for_check.scala 426:51:@457.4]
  assign _T_895 = stripe_cnt_inc == _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 426:51:@457.4]
  assign is_stripe_equal = is_batch_end & _T_895; // @[NV_NVDLA_CSC_dl_for_check.scala 426:33:@458.4]
  assign is_stripe_end = is_stripe_equal & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 427:34:@460.4]
  assign _T_898 = dat_exec_valid & is_batch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 428:52:@462.4]
  assign stripe_cnt_reg_en = layer_st | _T_898; // @[NV_NVDLA_CSC_dl_for_check.scala 428:34:@463.4]
  assign _T_900 = ~ is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 432:41:@465.6]
  assign _T_901 = is_stripe_equal & _T_900; // @[NV_NVDLA_CSC_dl_for_check.scala 432:39:@466.6]
  assign _T_903 = is_stripe_end ? 8'h0 : stripe_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 433:22:@467.6]
  assign _T_904 = _T_901 ? {{1'd0}, stripe_cnt} : _T_903; // @[NV_NVDLA_CSC_dl_for_check.scala 432:22:@468.6]
  assign _T_905 = layer_st ? 8'h0 : _T_904; // @[NV_NVDLA_CSC_dl_for_check.scala 431:22:@469.6]
  assign _GEN_66 = stripe_cnt_reg_en ? _T_905 : {{1'd0}, stripe_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 430:24:@464.4]
  assign dat_pipe_valid = dl_pvld | dat_pipe_local_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 446:27:@480.4]
  assign _T_914 = dat_pipe_valid & is_stripe_equal; // @[NV_NVDLA_CSC_dl_for_check.scala 443:49:@477.4]
  assign _T_917 = dl_pvld ? 1'h1 : dat_pipe_local_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 444:32:@478.4]
  assign dat_pipe_local_valid_w = _T_914 ? 1'h0 : _T_917; // @[NV_NVDLA_CSC_dl_for_check.scala 443:33:@479.4]
  assign dat_req_bytes = {1'h0,dl_channel_size}; // @[Cat.scala 30:58:@497.4]
  assign _GEN_67 = dat_exec_valid ? dat_req_bytes : dat_req_bytes_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 458:21:@498.4]
  assign _GEN_684 = {{10'd0}, sub_h_cmp_g1}; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@503.4]
  assign _T_941 = dataout_w_cnt + _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@503.4]
  assign dataout_w_cnt_inc = dataout_w_cnt + _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 468:39:@504.4]
  assign _T_942 = is_batch_end & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 469:29:@505.4]
  assign _T_943 = dataout_w_cnt >= dataout_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 469:61:@506.4]
  assign is_w_end = _T_942 & _T_943; // @[NV_NVDLA_CSC_dl_for_check.scala 469:44:@507.4]
  assign _T_945 = ~ dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 472:43:@510.4]
  assign _T_946 = is_stripe_end & _T_945; // @[NV_NVDLA_CSC_dl_for_check.scala 472:41:@511.4]
  assign _T_947 = is_w_end ? {{9'd0}, dataout_w_init} : dataout_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 473:26:@512.4]
  assign _T_948 = _T_946 ? dataout_w_ori : _T_947; // @[NV_NVDLA_CSC_dl_for_check.scala 472:26:@513.4]
  assign dataout_w_cnt_w = layer_st ? {{9'd0}, dataout_w_init} : _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 471:26:@514.4]
  assign _T_950 = _T_898 & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 474:70:@516.4]
  assign dataout_w_cnt_reg_en = layer_st | _T_950; // @[NV_NVDLA_CSC_dl_for_check.scala 474:37:@517.4]
  assign _T_951 = dat_exec_valid & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 475:55:@518.4]
  assign _T_952 = _T_951 & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 475:71:@519.4]
  assign dataout_w_ori_reg_en = layer_st | _T_952; // @[NV_NVDLA_CSC_dl_for_check.scala 475:37:@520.4]
  assign _GEN_68 = dataout_w_cnt_reg_en ? dataout_w_cnt_w : dataout_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 477:27:@521.4]
  assign _GEN_69 = dataout_w_ori_reg_en ? dataout_w_cnt_w : dataout_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 480:27:@524.4]
  assign is_last_channel = datain_c_cnt == datain_channel_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 487:37:@528.4]
  assign _T_956 = _T_951 & dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 488:70:@530.4]
  assign datain_c_cnt_reg_en = layer_st | _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 488:36:@531.4]
  assign _T_960 = datain_c_cnt + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@533.6]
  assign _T_961 = datain_c_cnt + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 493:34:@534.6]
  assign _T_962 = dl_channel_end ? 11'h0 : _T_961; // @[NV_NVDLA_CSC_dl_for_check.scala 492:24:@535.6]
  assign _T_963 = layer_st ? 11'h0 : _T_962; // @[NV_NVDLA_CSC_dl_for_check.scala 491:24:@536.6]
  assign _GEN_70 = datain_c_cnt_reg_en ? _T_963 : datain_c_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 490:26:@532.4]
  assign _GEN_685 = {{8'd0}, reg2dp_pad_left}; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@548.4]
  assign _T_983 = 13'h0 - _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@548.4]
  assign _T_984 = $unsigned(_T_983); // @[NV_NVDLA_CSC_dl_for_check.scala 508:41:@549.4]
  assign datain_w_cnt_st = is_img ? 14'h0 : _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 507:26:@550.4]
  assign _GEN_686 = {{10'd0}, conv_x_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@551.4]
  assign _T_985 = datain_w_cnt + _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@551.4]
  assign datain_w_cnt_inc = datain_w_cnt + _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 509:37:@552.4]
  assign _T_988 = is_w_end ? datain_w_cnt_st : datain_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 514:25:@555.4]
  assign _T_989 = _T_946 ? datain_w_ori : _T_988; // @[NV_NVDLA_CSC_dl_for_check.scala 513:25:@556.4]
  assign datain_w_cnt_w = layer_st ? datain_w_cnt_st : _T_989; // @[NV_NVDLA_CSC_dl_for_check.scala 512:25:@557.4]
  assign _GEN_687 = {{1'd0}, dl_w_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@558.4]
  assign dl_w_offset_ext = _GEN_687 * x_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 516:35:@558.4]
  assign _GEN_688 = {{3'd0}, dl_w_offset_ext}; // @[NV_NVDLA_CSC_dl_for_check.scala 517:34:@559.4]
  assign _T_990 = datain_w_cnt + _GEN_688; // @[NV_NVDLA_CSC_dl_for_check.scala 517:34:@559.4]
  assign datain_w_cur = _T_990[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 517:53:@560.4]
  assign _T_993 = is_img_d1[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 518:96:@563.4]
  assign _T_994 = ~ _T_993; // @[NV_NVDLA_CSC_dl_for_check.scala 518:86:@564.4]
  assign _T_995 = _T_950 & _T_994; // @[NV_NVDLA_CSC_dl_for_check.scala 518:84:@565.4]
  assign datain_w_cnt_reg_en = layer_st | _T_995; // @[NV_NVDLA_CSC_dl_for_check.scala 518:36:@566.4]
  assign _T_998 = is_img_d1[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 519:99:@569.4]
  assign _T_999 = ~ _T_998; // @[NV_NVDLA_CSC_dl_for_check.scala 519:89:@570.4]
  assign _T_1000 = _T_952 & _T_999; // @[NV_NVDLA_CSC_dl_for_check.scala 519:87:@571.4]
  assign datain_w_ori_reg_en = layer_st | _T_1000; // @[NV_NVDLA_CSC_dl_for_check.scala 519:36:@572.4]
  assign pixel_x_cnt_add = is_sub_h_end ? pixel_x_add : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 522:26:@573.4]
  assign _T_1004 = _T_371 == 6'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 524:79:@575.4]
  assign _T_1008 = _T_681 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@578.4]
  assign _T_1009 = _T_681 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 525:74:@579.4]
  assign total_channel_op = _T_1004 ? _T_681 : _T_1009; // @[NV_NVDLA_CSC_dl_for_check.scala 524:27:@580.4]
  assign _T_1010 = dl_channel_end & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 526:37:@581.4]
  assign _T_1012 = dl_block_end & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 527:35:@582.4]
  assign _T_1014 = channel_op_cnt + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 527:66:@583.4]
  assign _T_1015 = _T_1012 ? _T_1014 : {{1'd0}, channel_op_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 527:22:@584.4]
  assign _T_1016 = _T_1010 ? 14'h2 : _T_1015; // @[NV_NVDLA_CSC_dl_for_check.scala 526:22:@585.4]
  assign _GEN_689 = {{6'd0}, total_channel_op}; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@587.4]
  assign next_is_last_channel = channel_op_cnt >= _GEN_689; // @[NV_NVDLA_CSC_dl_for_check.scala 529:44:@587.4]
  assign _T_1017 = is_stripe_end & dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 533:39:@588.4]
  assign _T_1018 = _T_1017 & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 533:54:@589.4]
  assign _T_1019 = _T_1018 & is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 533:71:@590.4]
  assign _T_1022 = ~ is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 534:73:@593.4]
  assign _T_1023 = _T_1018 & _T_1022; // @[NV_NVDLA_CSC_dl_for_check.scala 534:71:@594.4]
  assign _GEN_690 = {{4'd0}, pixel_ch_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@595.4]
  assign _T_1024 = pixel_w_ch_ori + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 534:99:@595.4]
  assign _T_1026 = _T_1017 & next_is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 535:54:@597.4]
  assign _GEN_691 = {{9'd0}, pixel_x_init_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@598.4]
  assign _T_1027 = pixel_w_ori + _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 535:90:@598.4]
  assign _T_1029 = ~ next_is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 536:56:@600.4]
  assign _T_1030 = _T_1017 & _T_1029; // @[NV_NVDLA_CSC_dl_for_check.scala 536:54:@601.4]
  assign _T_1032 = pixel_w_ori + 16'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 536:91:@602.4]
  assign _T_1033 = ~ dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 537:41:@603.4]
  assign _T_1034 = is_stripe_end & _T_1033; // @[NV_NVDLA_CSC_dl_for_check.scala 537:39:@604.4]
  assign _GEN_692 = {{8'd0}, pixel_x_cnt_add}; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@605.4]
  assign _T_1035 = pixel_w_cnt + _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 537:81:@605.4]
  assign _T_1036 = _T_1034 ? {{1'd0}, pixel_w_ori} : _T_1035; // @[NV_NVDLA_CSC_dl_for_check.scala 537:24:@606.4]
  assign _T_1037 = _T_1030 ? _T_1032 : _T_1036; // @[NV_NVDLA_CSC_dl_for_check.scala 536:24:@607.4]
  assign _T_1038 = _T_1026 ? _T_1027 : _T_1037; // @[NV_NVDLA_CSC_dl_for_check.scala 535:24:@608.4]
  assign _T_1039 = _T_1023 ? _T_1024 : _T_1038; // @[NV_NVDLA_CSC_dl_for_check.scala 534:24:@609.4]
  assign _T_1040 = _T_1019 ? {{10'd0}, pixel_x_init} : _T_1039; // @[NV_NVDLA_CSC_dl_for_check.scala 533:24:@610.4]
  assign _T_1041 = layer_st_d1 ? {{10'd0}, pixel_x_init} : _T_1040; // @[NV_NVDLA_CSC_dl_for_check.scala 532:24:@611.4]
  assign pixel_w_cnt_w = _T_1041[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 537:105:@612.4]
  assign _T_1047 = pixel_w_cnt[15:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 539:68:@614.4]
  assign pixel_w_cur = {5'h0,_T_1047}; // @[Cat.scala 30:58:@615.4]
  assign _T_1056 = is_img_d1[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 542:68:@626.4]
  assign _T_1057 = dat_exec_valid & _T_1056; // @[NV_NVDLA_CSC_dl_for_check.scala 542:57:@627.4]
  assign _T_1058 = _T_1057 & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 542:72:@628.4]
  assign _T_1059 = _T_1058 & dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 542:88:@629.4]
  assign _T_1060 = _T_1059 & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 542:103:@630.4]
  assign pixel_ch_ori_reg_en = layer_st_d1 | _T_1060; // @[NV_NVDLA_CSC_dl_for_check.scala 542:39:@631.4]
  assign _T_1062 = _T_993 & dl_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 544:42:@633.4]
  assign _T_1065 = pixel_force_clr_d1 ? 1'h0 : pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 544:74:@634.4]
  assign pixel_force_fetch = _T_1062 ? 1'h1 : _T_1065; // @[NV_NVDLA_CSC_dl_for_check.scala 544:28:@635.4]
  assign _T_1067 = _T_993 & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 545:36:@637.4]
  assign _T_1068 = pixel_force_fetch | pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 545:72:@638.4]
  assign pixel_force_clr = _T_1067 & _T_1068; // @[NV_NVDLA_CSC_dl_for_check.scala 545:51:@639.4]
  assign _GEN_71 = datain_w_cnt_reg_en ? datain_w_cnt_w : datain_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@640.4]
  assign _GEN_72 = datain_w_cnt_reg_en ? pixel_w_cnt_w : pixel_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@640.4]
  assign _GEN_73 = datain_w_ori_reg_en ? datain_w_cnt_w : datain_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@644.4]
  assign _GEN_74 = datain_w_ori_reg_en ? pixel_w_cnt_w : pixel_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 551:26:@644.4]
  assign _GEN_75 = pixel_ch_ori_reg_en ? pixel_w_cnt_w : pixel_w_ch_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 555:26:@648.4]
  assign _GEN_693 = {{9'd0}, reg2dp_pad_top}; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@653.4]
  assign _T_1074 = 14'h0 - _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@653.4]
  assign _T_1075 = $unsigned(_T_1074); // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@654.4]
  assign datain_h_cnt_st = _T_1075[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 564:41:@655.4]
  assign _GEN_694 = {{10'd0}, conv_y_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@656.4]
  assign _T_1076 = datain_h_cnt + _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@656.4]
  assign datain_h_cnt_inc = datain_h_cnt + _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 565:37:@657.4]
  assign _T_1077 = is_stripe_end & dl_group_end; // @[NV_NVDLA_CSC_dl_for_check.scala 566:52:@658.4]
  assign _T_1078 = layer_st | _T_1077; // @[NV_NVDLA_CSC_dl_for_check.scala 566:35:@659.4]
  assign _T_1081 = is_w_end ? datain_h_cnt_inc : datain_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 568:25:@662.4]
  assign _T_1082 = _T_946 ? datain_h_ori : _T_1081; // @[NV_NVDLA_CSC_dl_for_check.scala 567:25:@663.4]
  assign datain_h_cnt_w = _T_1078 ? datain_h_cnt_st : _T_1082; // @[NV_NVDLA_CSC_dl_for_check.scala 566:25:@664.4]
  assign _T_1085 = _T_946 | is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 569:91:@667.4]
  assign _T_1086 = dat_exec_valid & _T_1085; // @[NV_NVDLA_CSC_dl_for_check.scala 569:54:@668.4]
  assign datain_h_cnt_reg_en = layer_st | _T_1086; // @[NV_NVDLA_CSC_dl_for_check.scala 569:36:@669.4]
  assign _GEN_695 = {{1'd0}, dl_h_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@673.4]
  assign dl_h_offset_ext = _GEN_695 * y_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 571:35:@673.4]
  assign _GEN_696 = {{3'd0}, dl_h_offset_ext}; // @[NV_NVDLA_CSC_dl_for_check.scala 572:34:@674.4]
  assign _T_1089 = datain_h_cnt + _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 572:34:@674.4]
  assign _GEN_697 = {{13'd0}, sub_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 572:53:@675.4]
  assign _T_1090 = _T_1089 + _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 572:53:@675.4]
  assign datain_h_cur = _T_1090[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 572:66:@676.4]
  assign _GEN_76 = datain_h_cnt_reg_en ? datain_h_cnt_w : datain_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 574:26:@677.4]
  assign _GEN_77 = dataout_w_ori_reg_en ? datain_h_cnt_w : datain_h_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 575:26:@680.4]
  assign _T_1091 = datain_w_cur[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 578:39:@683.4]
  assign _GEN_698 = {{1'd0}, datain_width_cmp}; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@684.4]
  assign _T_1092 = datain_w_cur > _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 578:59:@684.4]
  assign _T_1093 = _T_1091 | _T_1092; // @[NV_NVDLA_CSC_dl_for_check.scala 578:44:@685.4]
  assign _T_1094 = datain_h_cur[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 578:92:@686.4]
  assign _T_1095 = _T_1093 | _T_1094; // @[NV_NVDLA_CSC_dl_for_check.scala 578:78:@687.4]
  assign _GEN_699 = {{1'd0}, datain_height_cmp}; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@688.4]
  assign _T_1096 = datain_h_cur > _GEN_699; // @[NV_NVDLA_CSC_dl_for_check.scala 578:112:@688.4]
  assign dat_conv_req_dummy = _T_1095 | _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 578:97:@689.4]
  assign dat_img_req_dummy = _T_1094 | _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 581:42:@699.4]
  assign _T_1179 = is_img_d1[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 666:33:@785.4]
  assign _T_1180 = ~ is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 667:24:@786.4]
  assign _T_1182 = datain_w_cur[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 667:77:@787.4]
  assign _T_1183 = {2'h0,_T_1182}; // @[Cat.scala 30:58:@788.4]
  assign _T_1185 = dat_req_bytes > 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 668:38:@789.4]
  assign _T_1190 = datain_w_cur[12:1]; // @[NV_NVDLA_CSC_dl_for_check.scala 669:54:@792.4]
  assign _T_1191 = {3'h0,_T_1190}; // @[Cat.scala 30:58:@793.4]
  assign _T_1192 = _T_1185 ? _T_1183 : _T_1191; // @[NV_NVDLA_CSC_dl_for_check.scala 668:23:@794.4]
  assign _T_1193 = _T_1180 ? _T_1183 : _T_1192; // @[NV_NVDLA_CSC_dl_for_check.scala 667:23:@795.4]
  assign w_bias_int8 = _T_1179 ? pixel_w_cur : _T_1193; // @[NV_NVDLA_CSC_dl_for_check.scala 666:23:@796.4]
  assign w_bias_w = w_bias_int8[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 678:24:@798.4]
  assign _T_1108 = w_bias_w[13:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 585:32:@701.4]
  assign _GEN_701 = {{3'd0}, _T_1108}; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@702.4]
  assign dat_img_req_skip = _GEN_701 > entries_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 585:40:@702.4]
  assign _T_1109 = is_img_d1[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 586:34:@703.4]
  assign dat_req_dummy = _T_1109 ? dat_img_req_dummy : dat_conv_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 586:24:@704.4]
  assign _T_1110 = is_img_d1[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 587:29:@705.4]
  assign dat_req_skip = _T_1110 & dat_img_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 587:33:@706.4]
  assign _T_1111 = ~ dat_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 588:39:@707.4]
  assign _T_1112 = dat_exec_valid & _T_1111; // @[NV_NVDLA_CSC_dl_for_check.scala 588:37:@708.4]
  assign _T_1113 = ~ dat_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 588:56:@709.4]
  assign dat_req_valid = _T_1112 & _T_1113; // @[NV_NVDLA_CSC_dl_for_check.scala 588:54:@710.4]
  assign _T_1114 = is_img_d1[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 591:37:@711.4]
  assign _T_1115 = ~ _T_1114; // @[NV_NVDLA_CSC_dl_for_check.scala 591:27:@712.4]
  assign _T_1116 = datain_c_cnt[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 591:54:@713.4]
  assign dat_req_sub_c_w = _T_1115 ? _T_1116 : dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 591:26:@714.4]
  assign dat_req_sub_w_w = datain_w_cur[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 592:35:@715.4]
  assign _T_1118 = sub_h_cnt == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 593:55:@716.4]
  assign dat_req_sub_w_st_en = dat_exec_valid & _T_1118; // @[NV_NVDLA_CSC_dl_for_check.scala 593:42:@717.4]
  assign dat_req_stripe_end = is_stripe_equal & dat_pipe_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 596:42:@719.4]
  assign dat_req_flag_w = {dl_layer_end,dl_channel_end,dat_req_stripe_end,dl_pvld,batch_cnt}; // @[Cat.scala 30:58:@723.4]
  assign _T_1142 = dl_dat_release & is_stripe_equal; // @[NV_NVDLA_CSC_dl_for_check.scala 623:38:@743.6]
  assign _T_1143 = _T_1142 & dat_pipe_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 623:56:@744.6]
  assign _GEN_78 = dat_exec_valid ? dat_req_sub_w_w : dat_req_sub_w_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_79 = dat_exec_valid ? sub_h_cnt : dat_req_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_80 = dat_exec_valid ? dat_req_sub_c_w : dat_req_sub_c_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_81 = dat_exec_valid ? is_last_channel : dat_req_ch_end_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_82 = dat_exec_valid ? dat_exec_valid : dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_83 = dat_exec_valid ? dl_cur_sub_h : dat_req_cur_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_84 = dat_exec_valid ? dat_req_flag_w : {{1'd0}, dat_req_flag_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_85 = dat_exec_valid ? _T_1143 : dat_req_rls_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_86 = dat_exec_valid ? pixel_force_fetch : pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_87 = dat_exec_valid ? pixel_force_clr : pixel_force_clr_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 615:21:@735.4]
  assign _GEN_88 = dat_req_sub_w_st_en ? dl_pvld : dat_req_sub_w_st_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 627:26:@749.4]
  assign _T_1158 = is_img_d1[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 644:32:@759.4]
  assign _T_1159 = ~ _T_1158; // @[NV_NVDLA_CSC_dl_for_check.scala 644:22:@760.4]
  assign _T_1160 = datain_width[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 644:49:@761.4]
  assign c_bias_add = _T_1159 ? _T_1160 : 12'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 644:21:@762.4]
  assign _T_1163 = is_stripe_end & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 646:34:@763.4]
  assign _GEN_702 = {{1'd0}, c_bias_add}; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@764.4]
  assign _T_1165 = c_bias + _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@764.4]
  assign _T_1166 = c_bias + _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 646:64:@765.4]
  assign _T_1167 = _T_1163 ? 13'h0 : _T_1166; // @[NV_NVDLA_CSC_dl_for_check.scala 646:19:@766.4]
  assign c_bias_w = layer_st ? 13'h0 : _T_1167; // @[NV_NVDLA_CSC_dl_for_check.scala 645:19:@767.4]
  assign c_bias_d1_reg_en = c_bias != c_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 648:31:@771.4]
  assign _GEN_703 = {{2'd0}, h_bias_0_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@772.4]
  assign _T_1170 = datain_h_cnt * _GEN_703; // @[NV_NVDLA_CSC_dl_for_check.scala 651:32:@772.4]
  assign h_bias_0_w = _T_1170[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 651:50:@773.4]
  assign _GEN_704 = {{7'd0}, dl_h_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@774.4]
  assign _T_1171 = _GEN_704 * h_bias_1_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 652:31:@774.4]
  assign h_bias_1_w = _T_1171[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 652:49:@775.4]
  assign _GEN_705 = {{9'd0}, batch_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@776.4]
  assign _T_1172 = _GEN_705 * h_bias_2_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 653:29:@776.4]
  assign h_bias_2_w = _T_1172[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 653:47:@777.4]
  assign _T_1174 = _GEN_697 * h_bias_3_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 654:79:@778.4]
  assign _T_1175 = layer_st ? 17'h0 : _T_1174; // @[NV_NVDLA_CSC_dl_for_check.scala 654:21:@779.4]
  assign h_bias_3_w = _T_1175[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 654:97:@780.4]
  assign _T_1176 = is_img_d1[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 655:45:@781.4]
  assign _T_1177 = layer_st | _T_1176; // @[NV_NVDLA_CSC_dl_for_check.scala 655:34:@782.4]
  assign h_bias_reg_en = {_T_1177,dat_exec_valid}; // @[Cat.scala 30:58:@783.4]
  assign _GEN_89 = datain_c_cnt_reg_en ? c_bias_w : c_bias; // @[NV_NVDLA_CSC_dl_for_check.scala 682:20:@800.4]
  assign _GEN_90 = c_bias_d1_reg_en ? c_bias : c_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 685:23:@803.4]
  assign _T_1196 = h_bias_reg_en[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 688:19:@806.4]
  assign _GEN_91 = _T_1196 ? h_bias_0_w : h_bias_0_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@807.4]
  assign _GEN_92 = _T_1196 ? h_bias_1_w : h_bias_1_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@807.4]
  assign _GEN_93 = _T_1196 ? h_bias_2_w : h_bias_2_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@807.4]
  assign _T_1197 = h_bias_reg_en[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 693:19:@812.4]
  assign _GEN_94 = _T_1197 ? h_bias_3_w : h_bias_3_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 693:23:@813.4]
  assign _GEN_95 = dat_exec_valid ? w_bias_w : {{1'd0}, w_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 696:20:@816.4]
  assign _T_1288 = h_bias_0_d1 + h_bias_1_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 720:30:@844.4]
  assign _GEN_707 = {{1'd0}, h_bias_2_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 720:45:@845.4]
  assign _T_1289 = _T_1288 + _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 720:45:@845.4]
  assign _GEN_708 = {{2'd0}, h_bias_3_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 720:60:@846.4]
  assign _T_1290 = _T_1289 + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 720:60:@846.4]
  assign h_bias_d1 = _T_1290[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 720:75:@847.4]
  assign _GEN_709 = {{2'd0}, c_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@848.4]
  assign _T_1291 = dat_entry_st + _GEN_709; // @[NV_NVDLA_CSC_dl_for_check.scala 721:40:@848.4]
  assign _GEN_710 = {{3'd0}, h_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 721:53:@849.4]
  assign _T_1292 = _T_1291 + _GEN_710; // @[NV_NVDLA_CSC_dl_for_check.scala 721:53:@849.4]
  assign _GEN_711 = {{4'd0}, w_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 721:66:@850.4]
  assign dat_req_addr_sum = _T_1292 + _GEN_711; // @[NV_NVDLA_CSC_dl_for_check.scala 721:66:@850.4]
  assign _GEN_712 = {{4'd0}, _T_726}; // @[NV_NVDLA_CSC_dl_for_check.scala 722:45:@853.4]
  assign is_dat_req_addr_wrap = dat_req_addr_sum >= _GEN_712; // @[NV_NVDLA_CSC_dl_for_check.scala 722:45:@853.4]
  assign _T_1305 = dat_req_addr_sum - _GEN_712; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@856.4]
  assign _T_1306 = $unsigned(_T_1305); // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@857.4]
  assign dat_req_addr_wrap = _T_1306[17:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 723:42:@858.4]
  assign _T_1307 = layer_st | dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 724:35:@859.4]
  assign _T_1313 = dat_req_addr_sum[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 725:83:@861.4]
  assign _T_1314 = is_dat_req_addr_wrap ? dat_req_addr_wrap : {{5'd0}, _T_1313}; // @[NV_NVDLA_CSC_dl_for_check.scala 725:25:@862.4]
  assign dat_req_addr_w = _T_1307 ? 18'h1fff : _T_1314; // @[NV_NVDLA_CSC_dl_for_check.scala 724:25:@863.4]
  assign _T_1333 = 2'h2 == dat_req_sub_h_d1; // @[Mux.scala 46:19:@873.4]
  assign _T_1334 = _T_1333 ? dat_req_sub_h_addr_2 : 13'h0; // @[Mux.scala 46:16:@874.4]
  assign _T_1335 = 2'h1 == dat_req_sub_h_d1; // @[Mux.scala 46:19:@875.4]
  assign _T_1336 = _T_1335 ? dat_req_sub_h_addr_1 : _T_1334; // @[Mux.scala 46:16:@876.4]
  assign _T_1337 = 2'h0 == dat_req_sub_h_d1; // @[Mux.scala 46:19:@877.4]
  assign dat_req_addr_last = _T_1337 ? dat_req_sub_h_addr_0 : _T_1336; // @[Mux.scala 46:16:@878.4]
  assign _GEN_715 = {{5'd0}, dat_req_addr_last}; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@879.4]
  assign _T_1338 = _GEN_715 != dat_req_addr_w; // @[NV_NVDLA_CSC_dl_for_check.scala 732:65:@879.4]
  assign _T_1339 = _T_1338 | pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 732:85:@880.4]
  assign sc2buf_dat_rd_en_w = dat_req_valid_d1 & _T_1339; // @[NV_NVDLA_CSC_dl_for_check.scala 732:43:@881.4]
  assign _T_1340 = dat_req_valid_d1 | dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 734:38:@882.4]
  assign _T_1342 = dat_req_sub_h_d1 == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@883.4]
  assign _T_1343 = _T_1340 & _T_1342; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@884.4]
  assign dat_req_sub_h_addr_en_0 = layer_st | _T_1343; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@885.4]
  assign _T_1347 = dat_req_sub_h_d1 == 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@887.4]
  assign _T_1348 = _T_1340 & _T_1347; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@888.4]
  assign dat_req_sub_h_addr_en_1 = layer_st | _T_1348; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@889.4]
  assign _T_1352 = dat_req_sub_h_d1 == 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 734:78:@891.4]
  assign _T_1353 = _T_1340 & _T_1352; // @[NV_NVDLA_CSC_dl_for_check.scala 734:58:@892.4]
  assign dat_req_sub_h_addr_en_2 = layer_st | _T_1353; // @[NV_NVDLA_CSC_dl_for_check.scala 734:17:@893.4]
  assign _GEN_96 = dat_req_sub_h_addr_en_0 ? dat_req_addr_w : {{5'd0}, dat_req_sub_h_addr_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@903.4]
  assign _GEN_97 = dat_req_sub_h_addr_en_1 ? dat_req_addr_w : {{5'd0}, dat_req_sub_h_addr_1}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@906.4]
  assign _GEN_98 = dat_req_sub_h_addr_en_2 ? dat_req_addr_w : {{5'd0}, dat_req_sub_h_addr_2}; // @[NV_NVDLA_CSC_dl_for_check.scala 741:35:@909.4]
  assign _T_1369 = layer_st | sc2buf_dat_rd_en_w; // @[NV_NVDLA_CSC_dl_for_check.scala 747:14:@916.4]
  assign _GEN_100 = _T_1369 ? dat_req_addr_w : sc2buf_dat_rd_addr_out; // @[NV_NVDLA_CSC_dl_for_check.scala 747:34:@917.4]
  assign _GEN_101 = dat_exec_valid_d1 ? dat_req_sub_w_d1 : dat_req_pipe_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_102 = dat_exec_valid_d1 ? dat_req_sub_h_d1 : dat_req_pipe_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_103 = dat_exec_valid_d1 ? dat_req_sub_c_d1 : dat_req_pipe_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_104 = dat_exec_valid_d1 ? dat_req_ch_end_d1 : dat_req_pipe_ch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_105 = dat_exec_valid_d1 ? dat_req_bytes_d1 : dat_req_pipe_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_106 = dat_exec_valid_d1 ? dat_req_dummy_d1 : dat_req_pipe_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_107 = dat_exec_valid_d1 ? dat_req_cur_sub_h_d1 : dat_req_pipe_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_108 = dat_exec_valid_d1 ? dat_req_sub_w_st_d1 : dat_req_pipe_sub_w_st; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_109 = dat_exec_valid_d1 ? dat_req_rls_d1 : dat_req_pipe_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _GEN_110 = dat_exec_valid_d1 ? dat_req_flag_d1 : {{8'd0}, dat_exec_valid_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 754:24:@924.4]
  assign _T_1379 = {1'h0,dat_req_pipe_ch_end,dat_req_pipe_sub_c,dat_req_pipe_sub_h,dat_req_pipe_sub_w}; // @[Cat.scala 30:58:@944.4]
  assign dat_req_pipe_pd = {dat_req_pipe_flag,dat_req_pipe_rls,dat_req_pipe_sub_w_st,dat_req_pipe_dummy,dat_req_pipe_cur_sub_h,dat_req_pipe_bytes,_T_1379}; // @[Cat.scala 30:58:@950.4]
  assign _GEN_111 = dat_req_pipe_pvld ? dat_req_pipe_pd : _T_1408; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@992.4]
  assign _GEN_114 = _T_1389 ? _T_1408 : _T_1411; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1001.4]
  assign _GEN_117 = _T_1392 ? _T_1411 : _T_1414; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1010.4]
  assign _GEN_120 = _T_1395 ? _T_1414 : _T_1417; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1019.4]
  assign _GEN_123 = _T_1398 ? _T_1417 : _T_1420; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1028.4]
  assign _GEN_126 = _T_1401 ? _T_1420 : dat_rsp_pipe_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 799:33:@1037.4]
  assign dat_rsp_pipe_sub_w = dat_rsp_pipe_pd[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 816:41:@1045.4]
  assign dat_rsp_pipe_sub_h = dat_rsp_pipe_pd[3:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 817:41:@1046.4]
  assign dat_rsp_pipe_sub_c = dat_rsp_pipe_pd[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 818:41:@1047.4]
  assign dat_rsp_pipe_ch_end = dat_rsp_pipe_pd[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 819:42:@1048.4]
  assign dat_rsp_pipe_bytes = dat_rsp_pipe_pd[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 820:41:@1049.4]
  assign dat_rsp_pipe_cur_sub_h = dat_rsp_pipe_pd[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 821:45:@1050.4]
  assign dat_rsp_pipe_rls = dat_rsp_pipe_pd[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 824:39:@1053.4]
  assign dat_rsp_pipe_flag = dat_rsp_pipe_pd[28:20]; // @[NV_NVDLA_CSC_dl_for_check.scala 825:40:@1054.4]
  assign _T_1515 = is_img_d1[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 855:69:@1082.4]
  assign _T_1516 = _T_1515 & sc2buf_dat_rd_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 855:74:@1083.4]
  assign _T_1517 = ~ dat_l0c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 855:90:@1084.4]
  assign dat_l0c1_en = _T_1516 & _T_1517; // @[NV_NVDLA_CSC_dl_for_check.scala 855:88:@1085.4]
  assign _T_1546 = sc2buf_dat_rd_valid ? 1'h0 : dat_l0c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 870:22:@1119.4]
  assign _T_1560 = sc2buf_dat_rd_valid ? dat_l0c0_dummy : dat_l0c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 874:48:@1130.4]
  assign _T_1561 = dat_l0c1_en ? 1'h0 : _T_1560; // @[NV_NVDLA_CSC_dl_for_check.scala 874:22:@1131.4]
  assign _T_1626 = {dat_rsp_pipe_flag,dat_rsp_pipe_rls,dat_rsp_pipe_cur_sub_h,dat_rsp_pipe_bytes,1'h0,dat_rsp_pipe_ch_end,dat_rsp_pipe_sub_c,dat_rsp_pipe_sub_h,dat_rsp_pipe_sub_w}; // @[Cat.scala 30:58:@1198.4]
  assign _GEN_137 = dat_rsp_pipe_pvld ? _T_1626 : _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1201.4]
  assign _GEN_138 = dat_rsp_l0_pvld ? _T_1608 : _T_1611; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1205.4]
  assign _GEN_139 = dat_rsp_l1_pvld ? _T_1611 : _T_1614; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1209.4]
  assign _GEN_140 = dat_rsp_l2_pvld ? _T_1614 : _T_1617; // @[NV_NVDLA_CSC_dl_for_check.scala 913:28:@1213.4]
  assign dat_rsp_l0_sub_c = _T_1608[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 931:39:@1239.4]
  assign dat_rsp_l1_sub_c = _T_1611[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 932:39:@1240.4]
  assign dat_rsp_l2_sub_c = _T_1614[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 933:39:@1241.4]
  assign dat_rsp_l3_sub_c = _T_1617[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 934:39:@1242.4]
  assign dat_rsp_l0_flag = _T_1608[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 936:38:@1243.4]
  assign dat_rsp_l1_flag = _T_1611[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 937:38:@1244.4]
  assign dat_rsp_l2_flag = _T_1614[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 938:38:@1245.4]
  assign dat_rsp_l3_flag = _T_1617[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 939:38:@1246.4]
  assign dat_rsp_l0_stripe_end = dat_rsp_l0_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 941:44:@1247.4]
  assign dat_rsp_l1_stripe_end = dat_rsp_l1_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 942:44:@1248.4]
  assign dat_rsp_l2_stripe_end = dat_rsp_l2_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 943:44:@1249.4]
  assign dat_rsp_l3_stripe_end = dat_rsp_l3_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 944:44:@1250.4]
  assign dat_rsp_sub_w = dat_rsp_pd[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 947:31:@1251.4]
  assign dat_rsp_bytes = dat_rsp_pd[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 951:31:@1255.4]
  assign dat_rsp_cur_sub_h = dat_rsp_pd[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 952:35:@1256.4]
  assign dat_rsp_flag = dat_rsp_pd[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 954:30:@1259.4]
  assign rsp_sft_cnt_l0_sub = sc2buf_dat_rd_valid ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 963:29:@1265.4]
  assign _T_1664 = pixel_x_byte_stride > 7'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 968:50:@1269.4]
  assign _GEN_716 = {{1'd0}, pixel_x_byte_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1270.4]
  assign _T_1666 = rsp_sft_cnt_l0 + _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 968:111:@1270.4]
  assign _GEN_717 = {{1'd0}, rsp_sft_cnt_l0_sub}; // @[NV_NVDLA_CSC_dl_for_check.scala 968:134:@1271.4]
  assign _T_1667 = _T_1666 - _GEN_717; // @[NV_NVDLA_CSC_dl_for_check.scala 968:134:@1271.4]
  assign _T_1668 = $unsigned(_T_1667); // @[NV_NVDLA_CSC_dl_for_check.scala 968:134:@1272.4]
  assign _T_1669 = _T_1664 ? 10'h40 : _T_1668; // @[NV_NVDLA_CSC_dl_for_check.scala 968:29:@1273.4]
  assign rsp_sft_cnt_l0_inc = _T_1669[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 968:156:@1274.4]
  assign _T_1673 = rsp_sft_cnt_l1 + _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 969:111:@1276.4]
  assign _T_1674 = _T_1673 - 9'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 969:134:@1277.4]
  assign _T_1675 = $unsigned(_T_1674); // @[NV_NVDLA_CSC_dl_for_check.scala 969:134:@1278.4]
  assign _T_1676 = _T_1664 ? 10'h40 : _T_1675; // @[NV_NVDLA_CSC_dl_for_check.scala 969:29:@1279.4]
  assign rsp_sft_cnt_l1_inc = _T_1676[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 969:156:@1280.4]
  assign _T_1680 = rsp_sft_cnt_l2 + _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 970:111:@1282.4]
  assign _T_1681 = {{1'd0}, _T_1680}; // @[NV_NVDLA_CSC_dl_for_check.scala 970:134:@1283.4]
  assign _T_1682 = _T_1664 ? 10'h40 : _T_1681; // @[NV_NVDLA_CSC_dl_for_check.scala 970:29:@1284.4]
  assign rsp_sft_cnt_l2_inc = _T_1682[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 970:156:@1285.4]
  assign _T_1686 = rsp_sft_cnt_l3 + _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 971:111:@1287.4]
  assign _T_1687 = {{1'd0}, _T_1686}; // @[NV_NVDLA_CSC_dl_for_check.scala 971:134:@1288.4]
  assign _T_1688 = _T_1664 ? 10'h40 : _T_1687; // @[NV_NVDLA_CSC_dl_for_check.scala 971:29:@1289.4]
  assign rsp_sft_cnt_l3_inc = _T_1688[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 971:156:@1290.4]
  assign _T_1690 = ~ dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 980:52:@1291.4]
  assign _T_1691 = dat_rsp_l0_stripe_end & _T_1690; // @[NV_NVDLA_CSC_dl_for_check.scala 980:50:@1292.4]
  assign _T_1692 = dat_rsp_l0_stripe_end & dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 981:50:@1293.4]
  assign _T_1697 = _T_1692 ? 8'h40 : rsp_sft_cnt_l0_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 981:27:@1296.4]
  assign _T_1698 = _T_1691 ? rsp_sft_cnt_l0_ori : _T_1697; // @[NV_NVDLA_CSC_dl_for_check.scala 980:27:@1297.4]
  assign rsp_sft_cnt_l0_w = layer_st ? 8'h40 : _T_1698; // @[NV_NVDLA_CSC_dl_for_check.scala 979:27:@1298.4]
  assign _T_1700 = ~ dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 985:52:@1299.4]
  assign _T_1701 = dat_rsp_l1_stripe_end & _T_1700; // @[NV_NVDLA_CSC_dl_for_check.scala 985:50:@1300.4]
  assign _T_1702 = dat_rsp_l1_stripe_end & dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 986:50:@1301.4]
  assign _T_1707 = _T_1702 ? 8'h40 : rsp_sft_cnt_l1_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 986:27:@1304.4]
  assign _T_1708 = _T_1701 ? rsp_sft_cnt_l1_ori : _T_1707; // @[NV_NVDLA_CSC_dl_for_check.scala 985:27:@1305.4]
  assign rsp_sft_cnt_l1_w = layer_st ? 8'h40 : _T_1708; // @[NV_NVDLA_CSC_dl_for_check.scala 984:27:@1306.4]
  assign _T_1710 = ~ dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 990:52:@1307.4]
  assign _T_1711 = dat_rsp_l2_stripe_end & _T_1710; // @[NV_NVDLA_CSC_dl_for_check.scala 990:50:@1308.4]
  assign _T_1712 = dat_rsp_l2_stripe_end & dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 991:50:@1309.4]
  assign _T_1717 = _T_1712 ? 8'h40 : rsp_sft_cnt_l2_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 991:27:@1312.4]
  assign _T_1718 = _T_1711 ? rsp_sft_cnt_l2_ori : _T_1717; // @[NV_NVDLA_CSC_dl_for_check.scala 990:27:@1313.4]
  assign rsp_sft_cnt_l2_w = layer_st ? 8'h40 : _T_1718; // @[NV_NVDLA_CSC_dl_for_check.scala 989:27:@1314.4]
  assign _T_1720 = ~ dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 995:52:@1315.4]
  assign _T_1721 = dat_rsp_l3_stripe_end & _T_1720; // @[NV_NVDLA_CSC_dl_for_check.scala 995:50:@1316.4]
  assign _T_1722 = dat_rsp_l3_stripe_end & dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 996:50:@1317.4]
  assign _T_1727 = _T_1722 ? 8'h40 : rsp_sft_cnt_l3_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 996:27:@1320.4]
  assign _T_1728 = _T_1721 ? rsp_sft_cnt_l3_ori : _T_1727; // @[NV_NVDLA_CSC_dl_for_check.scala 995:27:@1321.4]
  assign rsp_sft_cnt_l3_w = layer_st ? 8'h40 : _T_1728; // @[NV_NVDLA_CSC_dl_for_check.scala 994:27:@1322.4]
  assign _T_1729 = is_img_d1[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:46:@1323.4]
  assign _T_1730 = _T_1729 & dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:51:@1324.4]
  assign rsp_sft_cnt_l0_en = layer_st | _T_1730; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:34:@1325.4]
  assign _T_1731 = is_img_d1[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:46:@1326.4]
  assign _T_1732 = _T_1731 & dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:51:@1327.4]
  assign _T_1734 = sub_h_total_g5 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:87:@1328.4]
  assign _T_1735 = _T_1732 & _T_1734; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:69:@1329.4]
  assign rsp_sft_cnt_l1_en = layer_st | _T_1735; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:34:@1330.4]
  assign _T_1736 = is_img_d1[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:46:@1331.4]
  assign _T_1737 = _T_1736 & dat_rsp_l2_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:51:@1332.4]
  assign _T_1739 = sub_h_total_g5 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:87:@1333.4]
  assign _T_1740 = _T_1737 & _T_1739; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:69:@1334.4]
  assign rsp_sft_cnt_l2_en = layer_st | _T_1740; // @[NV_NVDLA_CSC_dl_for_check.scala 1002:34:@1335.4]
  assign _T_1741 = is_img_d1[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:46:@1336.4]
  assign _T_1742 = _T_1741 & dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:51:@1337.4]
  assign _T_1745 = _T_1742 & _T_1739; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:69:@1339.4]
  assign rsp_sft_cnt_l3_en = layer_st | _T_1745; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:34:@1340.4]
  assign _T_1746 = is_img_d1[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:50:@1341.4]
  assign _T_1747 = _T_1746 & dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:55:@1342.4]
  assign _T_1748 = _T_1747 & dat_rsp_l0_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:73:@1343.4]
  assign _T_1749 = _T_1748 & dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:97:@1344.4]
  assign rsp_sft_cnt_l0_ori_en = layer_st | _T_1749; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:38:@1345.4]
  assign _T_1750 = is_img_d1[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:50:@1346.4]
  assign _T_1751 = _T_1750 & dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:55:@1347.4]
  assign _T_1752 = _T_1751 & dat_rsp_l1_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:73:@1348.4]
  assign _T_1753 = _T_1752 & dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:97:@1349.4]
  assign _T_1755 = sub_h_total_g6 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:138:@1350.4]
  assign _T_1756 = _T_1753 & _T_1755; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:120:@1351.4]
  assign rsp_sft_cnt_l1_ori_en = layer_st | _T_1756; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:38:@1352.4]
  assign _T_1757 = is_img_d1[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:50:@1353.4]
  assign _T_1758 = _T_1757 & dat_rsp_l2_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:55:@1354.4]
  assign _T_1759 = _T_1758 & dat_rsp_l2_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:73:@1355.4]
  assign _T_1760 = _T_1759 & dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:97:@1356.4]
  assign _T_1762 = sub_h_total_g6 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:138:@1357.4]
  assign _T_1763 = _T_1760 & _T_1762; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:120:@1358.4]
  assign rsp_sft_cnt_l2_ori_en = layer_st | _T_1763; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:38:@1359.4]
  assign _T_1764 = is_img_d1[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:50:@1360.4]
  assign _T_1765 = _T_1764 & dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:55:@1361.4]
  assign _T_1766 = _T_1765 & dat_rsp_l3_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:73:@1362.4]
  assign _T_1767 = _T_1766 & dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:97:@1363.4]
  assign _T_1770 = _T_1767 & _T_1762; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:120:@1365.4]
  assign rsp_sft_cnt_l3_ori_en = layer_st | _T_1770; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:38:@1366.4]
  assign _GEN_141 = rsp_sft_cnt_l0_en ? rsp_sft_cnt_l0_w : rsp_sft_cnt_l0; // @[NV_NVDLA_CSC_dl_for_check.scala 1010:24:@1367.4]
  assign _GEN_142 = rsp_sft_cnt_l1_en ? rsp_sft_cnt_l1_w : rsp_sft_cnt_l1; // @[NV_NVDLA_CSC_dl_for_check.scala 1011:24:@1370.4]
  assign _GEN_143 = rsp_sft_cnt_l2_en ? rsp_sft_cnt_l2_w : rsp_sft_cnt_l2; // @[NV_NVDLA_CSC_dl_for_check.scala 1012:24:@1373.4]
  assign _GEN_144 = rsp_sft_cnt_l3_en ? rsp_sft_cnt_l3_w : rsp_sft_cnt_l3; // @[NV_NVDLA_CSC_dl_for_check.scala 1013:24:@1376.4]
  assign _GEN_145 = rsp_sft_cnt_l0_ori_en ? rsp_sft_cnt_l0_w : rsp_sft_cnt_l0_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1014:28:@1379.4]
  assign _GEN_146 = rsp_sft_cnt_l1_ori_en ? rsp_sft_cnt_l1_w : rsp_sft_cnt_l1_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1015:28:@1382.4]
  assign _GEN_147 = rsp_sft_cnt_l2_ori_en ? rsp_sft_cnt_l2_w : rsp_sft_cnt_l2_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1016:28:@1385.4]
  assign _GEN_148 = rsp_sft_cnt_l3_ori_en ? rsp_sft_cnt_l3_w : rsp_sft_cnt_l3_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1017:28:@1388.4]
  assign _T_1771 = pad_value[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:55:@1391.4]
  assign _T_1774 = {_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771}; // @[Cat.scala 30:58:@1394.4]
  assign _T_1775 = {_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1774}; // @[Cat.scala 30:58:@1395.4]
  assign _T_1776 = {_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1771,_T_1774,_T_1775}; // @[Cat.scala 30:58:@1396.4]
  assign dat_rsp_pad_value = {_T_1776,_T_1776}; // @[Cat.scala 30:58:@1397.4]
  assign dat_rsp_l0c0 = dat_l0c0_dummy ? dat_rsp_pad_value : dat_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1028:23:@1398.4]
  assign dat_rsp_l0c1 = dat_l0c1_dummy ? dat_rsp_pad_value : dat_l0c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1033:23:@1402.4]
  assign _T_1778 = is_img_d1[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:37:@1407.4]
  assign _T_1781 = dat_rsp_bytes <= 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:43:@1408.4]
  assign _T_1782 = dat_rsp_sub_w[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:87:@1409.4]
  assign _T_1784 = _T_1782 == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:91:@1410.4]
  assign _T_1785 = _T_1781 & _T_1784; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:72:@1411.4]
  assign _T_1787 = dat_rsp_l0c0[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:171:@1412.4]
  assign _T_1788 = {256'h0,_T_1787}; // @[Cat.scala 30:58:@1413.4]
  assign _T_1794 = _T_1781 & _T_1782; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:72:@1417.4]
  assign _T_1796 = dat_rsp_l0c0[511:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:171:@1418.4]
  assign _T_1797 = {256'h0,_T_1796}; // @[Cat.scala 30:58:@1419.4]
  assign _T_1798 = _T_1794 ? _T_1797 : dat_rsp_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1048:27:@1420.4]
  assign _T_1799 = _T_1785 ? _T_1788 : _T_1798; // @[NV_NVDLA_CSC_dl_for_check.scala 1047:27:@1421.4]
  assign dat_rsp_conv_8b = _T_1778 ? 512'h0 : _T_1799; // @[NV_NVDLA_CSC_dl_for_check.scala 1046:27:@1422.4]
  assign dat_rsp_conv_0 = dat_rsp_conv_8b[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1425.4]
  assign dat_rsp_conv_1 = dat_rsp_conv_8b[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1427.4]
  assign dat_rsp_conv_2 = dat_rsp_conv_8b[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1429.4]
  assign dat_rsp_conv_3 = dat_rsp_conv_8b[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1431.4]
  assign dat_rsp_conv_4 = dat_rsp_conv_8b[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1433.4]
  assign dat_rsp_conv_5 = dat_rsp_conv_8b[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1435.4]
  assign dat_rsp_conv_6 = dat_rsp_conv_8b[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1437.4]
  assign dat_rsp_conv_7 = dat_rsp_conv_8b[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1439.4]
  assign dat_rsp_conv_8 = dat_rsp_conv_8b[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1441.4]
  assign dat_rsp_conv_9 = dat_rsp_conv_8b[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1443.4]
  assign dat_rsp_conv_10 = dat_rsp_conv_8b[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1445.4]
  assign dat_rsp_conv_11 = dat_rsp_conv_8b[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1447.4]
  assign dat_rsp_conv_12 = dat_rsp_conv_8b[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1449.4]
  assign dat_rsp_conv_13 = dat_rsp_conv_8b[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1451.4]
  assign dat_rsp_conv_14 = dat_rsp_conv_8b[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1453.4]
  assign dat_rsp_conv_15 = dat_rsp_conv_8b[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1455.4]
  assign dat_rsp_conv_16 = dat_rsp_conv_8b[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1457.4]
  assign dat_rsp_conv_17 = dat_rsp_conv_8b[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1459.4]
  assign dat_rsp_conv_18 = dat_rsp_conv_8b[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1461.4]
  assign dat_rsp_conv_19 = dat_rsp_conv_8b[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1463.4]
  assign dat_rsp_conv_20 = dat_rsp_conv_8b[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1465.4]
  assign dat_rsp_conv_21 = dat_rsp_conv_8b[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1467.4]
  assign dat_rsp_conv_22 = dat_rsp_conv_8b[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1469.4]
  assign dat_rsp_conv_23 = dat_rsp_conv_8b[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1471.4]
  assign dat_rsp_conv_24 = dat_rsp_conv_8b[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1473.4]
  assign dat_rsp_conv_25 = dat_rsp_conv_8b[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1475.4]
  assign dat_rsp_conv_26 = dat_rsp_conv_8b[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1477.4]
  assign dat_rsp_conv_27 = dat_rsp_conv_8b[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1479.4]
  assign dat_rsp_conv_28 = dat_rsp_conv_8b[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1481.4]
  assign dat_rsp_conv_29 = dat_rsp_conv_8b[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1483.4]
  assign dat_rsp_conv_30 = dat_rsp_conv_8b[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1485.4]
  assign dat_rsp_conv_31 = dat_rsp_conv_8b[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1487.4]
  assign dat_rsp_conv_32 = dat_rsp_conv_8b[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1489.4]
  assign dat_rsp_conv_33 = dat_rsp_conv_8b[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1491.4]
  assign dat_rsp_conv_34 = dat_rsp_conv_8b[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1493.4]
  assign dat_rsp_conv_35 = dat_rsp_conv_8b[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1495.4]
  assign dat_rsp_conv_36 = dat_rsp_conv_8b[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1497.4]
  assign dat_rsp_conv_37 = dat_rsp_conv_8b[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1499.4]
  assign dat_rsp_conv_38 = dat_rsp_conv_8b[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1501.4]
  assign dat_rsp_conv_39 = dat_rsp_conv_8b[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1503.4]
  assign dat_rsp_conv_40 = dat_rsp_conv_8b[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1505.4]
  assign dat_rsp_conv_41 = dat_rsp_conv_8b[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1507.4]
  assign dat_rsp_conv_42 = dat_rsp_conv_8b[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1509.4]
  assign dat_rsp_conv_43 = dat_rsp_conv_8b[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1511.4]
  assign dat_rsp_conv_44 = dat_rsp_conv_8b[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1513.4]
  assign dat_rsp_conv_45 = dat_rsp_conv_8b[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1515.4]
  assign dat_rsp_conv_46 = dat_rsp_conv_8b[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1517.4]
  assign dat_rsp_conv_47 = dat_rsp_conv_8b[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1519.4]
  assign dat_rsp_conv_48 = dat_rsp_conv_8b[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1521.4]
  assign dat_rsp_conv_49 = dat_rsp_conv_8b[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1523.4]
  assign dat_rsp_conv_50 = dat_rsp_conv_8b[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1525.4]
  assign dat_rsp_conv_51 = dat_rsp_conv_8b[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1527.4]
  assign dat_rsp_conv_52 = dat_rsp_conv_8b[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1529.4]
  assign dat_rsp_conv_53 = dat_rsp_conv_8b[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1531.4]
  assign dat_rsp_conv_54 = dat_rsp_conv_8b[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1533.4]
  assign dat_rsp_conv_55 = dat_rsp_conv_8b[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1535.4]
  assign dat_rsp_conv_56 = dat_rsp_conv_8b[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1537.4]
  assign dat_rsp_conv_57 = dat_rsp_conv_8b[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1539.4]
  assign dat_rsp_conv_58 = dat_rsp_conv_8b[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1541.4]
  assign dat_rsp_conv_59 = dat_rsp_conv_8b[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1543.4]
  assign dat_rsp_conv_60 = dat_rsp_conv_8b[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1545.4]
  assign dat_rsp_conv_61 = dat_rsp_conv_8b[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1547.4]
  assign dat_rsp_conv_62 = dat_rsp_conv_8b[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1549.4]
  assign dat_rsp_conv_63 = dat_rsp_conv_8b[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1064:39:@1551.4]
  assign _T_1940 = is_img_d1[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:39:@1559.4]
  assign _T_1941 = ~ _T_1940; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:29:@1560.4]
  assign _T_1943 = {dat_rsp_l0c0,dat_rsp_l0c1}; // @[Cat.scala 30:58:@1561.4]
  assign dat_rsp_l0_sft_in = _T_1941 ? 1024'h0 : _T_1943; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:28:@1562.4]
  assign _T_1944 = is_img_d1[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:39:@1563.4]
  assign _T_1945 = ~ _T_1944; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:29:@1564.4]
  assign _T_1947 = {_T_1776,_T_1776,_T_1776,_T_1776}; // @[Cat.scala 30:58:@1565.4]
  assign dat_rsp_l1_sft_in = _T_1945 ? 1024'h0 : _T_1947; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:28:@1566.4]
  assign _T_1948 = is_img_d1[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:39:@1567.4]
  assign _T_1949 = ~ _T_1948; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:29:@1568.4]
  assign dat_rsp_l2_sft_in = _T_1949 ? 1024'h0 : _T_1947; // @[NV_NVDLA_CSC_dl_for_check.scala 1079:28:@1570.4]
  assign _T_1952 = is_img_d1[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:39:@1571.4]
  assign _T_1953 = ~ _T_1952; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:29:@1572.4]
  assign dat_rsp_l3_sft_in = _T_1953 ? 1024'h0 : _T_1947; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:28:@1574.4]
  assign _T_1957 = {rsp_sft_cnt_l0,3'h0}; // @[Cat.scala 30:58:@1575.4]
  assign _T_1958 = dat_rsp_l0_sft_in >> _T_1957; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:41:@1576.4]
  assign dat_rsp_l0_sft = _T_1958[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:82:@1577.4]
  assign _T_1960 = {rsp_sft_cnt_l1,3'h0}; // @[Cat.scala 30:58:@1578.4]
  assign _T_1961 = dat_rsp_l1_sft_in >> _T_1960; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:41:@1579.4]
  assign dat_rsp_l1_sft = _T_1961[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1083:82:@1580.4]
  assign _T_1963 = {rsp_sft_cnt_l2,3'h0}; // @[Cat.scala 30:58:@1581.4]
  assign _T_1964 = dat_rsp_l2_sft_in >> _T_1963; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:41:@1582.4]
  assign dat_rsp_l2_sft = _T_1964[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1084:82:@1583.4]
  assign _T_1966 = {rsp_sft_cnt_l3,3'h0}; // @[Cat.scala 30:58:@1584.4]
  assign _T_1967 = dat_rsp_l3_sft_in >> _T_1966; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:41:@1585.4]
  assign dat_rsp_l3_sft = _T_1967[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1085:82:@1586.4]
  assign _T_1968 = is_img_d1[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:36:@1587.4]
  assign _T_1969 = ~ _T_1968; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:26:@1588.4]
  assign _T_1972 = sub_h_total_g8 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:41:@1589.4]
  assign _T_1973 = dat_rsp_l3_sft[127:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:81:@1590.4]
  assign _T_1979 = {_T_1973,dat_rsp_l2_sft_d3,dat_rsp_l1_sft_d3,dat_rsp_l0_sft_d3}; // @[Cat.scala 30:58:@1596.4]
  assign _T_1981 = sub_h_total_g8 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:41:@1597.4]
  assign _T_1982 = dat_rsp_l1_sft[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:81:@1598.4]
  assign _T_1984 = {_T_1982,dat_rsp_l0_sft_d1}; // @[Cat.scala 30:58:@1600.4]
  assign _T_1986 = _T_1981 ? _T_1984 : dat_rsp_l0_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1089:25:@1602.4]
  assign _T_1987 = _T_1972 ? _T_1979 : _T_1986; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:25:@1603.4]
  assign dat_rsp_img_8b = _T_1969 ? 512'h0 : _T_1987; // @[NV_NVDLA_CSC_dl_for_check.scala 1087:25:@1604.4]
  assign dat_rsp_img_0 = dat_rsp_img_8b[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1606.4]
  assign dat_rsp_img_1 = dat_rsp_img_8b[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1608.4]
  assign dat_rsp_img_2 = dat_rsp_img_8b[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1610.4]
  assign dat_rsp_img_3 = dat_rsp_img_8b[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1612.4]
  assign dat_rsp_img_4 = dat_rsp_img_8b[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1614.4]
  assign dat_rsp_img_5 = dat_rsp_img_8b[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1616.4]
  assign dat_rsp_img_6 = dat_rsp_img_8b[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1618.4]
  assign dat_rsp_img_7 = dat_rsp_img_8b[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1620.4]
  assign dat_rsp_img_8 = dat_rsp_img_8b[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1622.4]
  assign dat_rsp_img_9 = dat_rsp_img_8b[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1624.4]
  assign dat_rsp_img_10 = dat_rsp_img_8b[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1626.4]
  assign dat_rsp_img_11 = dat_rsp_img_8b[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1628.4]
  assign dat_rsp_img_12 = dat_rsp_img_8b[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1630.4]
  assign dat_rsp_img_13 = dat_rsp_img_8b[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1632.4]
  assign dat_rsp_img_14 = dat_rsp_img_8b[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1634.4]
  assign dat_rsp_img_15 = dat_rsp_img_8b[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1636.4]
  assign dat_rsp_img_16 = dat_rsp_img_8b[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1638.4]
  assign dat_rsp_img_17 = dat_rsp_img_8b[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1640.4]
  assign dat_rsp_img_18 = dat_rsp_img_8b[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1642.4]
  assign dat_rsp_img_19 = dat_rsp_img_8b[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1644.4]
  assign dat_rsp_img_20 = dat_rsp_img_8b[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1646.4]
  assign dat_rsp_img_21 = dat_rsp_img_8b[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1648.4]
  assign dat_rsp_img_22 = dat_rsp_img_8b[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1650.4]
  assign dat_rsp_img_23 = dat_rsp_img_8b[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1652.4]
  assign dat_rsp_img_24 = dat_rsp_img_8b[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1654.4]
  assign dat_rsp_img_25 = dat_rsp_img_8b[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1656.4]
  assign dat_rsp_img_26 = dat_rsp_img_8b[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1658.4]
  assign dat_rsp_img_27 = dat_rsp_img_8b[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1660.4]
  assign dat_rsp_img_28 = dat_rsp_img_8b[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1662.4]
  assign dat_rsp_img_29 = dat_rsp_img_8b[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1664.4]
  assign dat_rsp_img_30 = dat_rsp_img_8b[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1666.4]
  assign dat_rsp_img_31 = dat_rsp_img_8b[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1668.4]
  assign dat_rsp_img_32 = dat_rsp_img_8b[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1670.4]
  assign dat_rsp_img_33 = dat_rsp_img_8b[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1672.4]
  assign dat_rsp_img_34 = dat_rsp_img_8b[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1674.4]
  assign dat_rsp_img_35 = dat_rsp_img_8b[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1676.4]
  assign dat_rsp_img_36 = dat_rsp_img_8b[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1678.4]
  assign dat_rsp_img_37 = dat_rsp_img_8b[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1680.4]
  assign dat_rsp_img_38 = dat_rsp_img_8b[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1682.4]
  assign dat_rsp_img_39 = dat_rsp_img_8b[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1684.4]
  assign dat_rsp_img_40 = dat_rsp_img_8b[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1686.4]
  assign dat_rsp_img_41 = dat_rsp_img_8b[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1688.4]
  assign dat_rsp_img_42 = dat_rsp_img_8b[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1690.4]
  assign dat_rsp_img_43 = dat_rsp_img_8b[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1692.4]
  assign dat_rsp_img_44 = dat_rsp_img_8b[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1694.4]
  assign dat_rsp_img_45 = dat_rsp_img_8b[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1696.4]
  assign dat_rsp_img_46 = dat_rsp_img_8b[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1698.4]
  assign dat_rsp_img_47 = dat_rsp_img_8b[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1700.4]
  assign dat_rsp_img_48 = dat_rsp_img_8b[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1702.4]
  assign dat_rsp_img_49 = dat_rsp_img_8b[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1704.4]
  assign dat_rsp_img_50 = dat_rsp_img_8b[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1706.4]
  assign dat_rsp_img_51 = dat_rsp_img_8b[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1708.4]
  assign dat_rsp_img_52 = dat_rsp_img_8b[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1710.4]
  assign dat_rsp_img_53 = dat_rsp_img_8b[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1712.4]
  assign dat_rsp_img_54 = dat_rsp_img_8b[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1714.4]
  assign dat_rsp_img_55 = dat_rsp_img_8b[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1716.4]
  assign dat_rsp_img_56 = dat_rsp_img_8b[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1718.4]
  assign dat_rsp_img_57 = dat_rsp_img_8b[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1720.4]
  assign dat_rsp_img_58 = dat_rsp_img_8b[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1722.4]
  assign dat_rsp_img_59 = dat_rsp_img_8b[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1724.4]
  assign dat_rsp_img_60 = dat_rsp_img_8b[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1726.4]
  assign dat_rsp_img_61 = dat_rsp_img_8b[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1728.4]
  assign dat_rsp_img_62 = dat_rsp_img_8b[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1730.4]
  assign dat_rsp_img_63 = dat_rsp_img_8b[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:37:@1732.4]
  assign _T_2122 = sub_h_total_g9 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:59:@1734.4]
  assign dat_rsp_sft_d1_en = dat_rsp_l0_pvld & _T_2122; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:41:@1735.4]
  assign _T_2124 = sub_h_total_g9 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:59:@1736.4]
  assign dat_rsp_sft_d2_en = dat_rsp_l1_pvld & _T_2124; // @[NV_NVDLA_CSC_dl_for_check.scala 1099:41:@1737.4]
  assign dat_rsp_sft_d3_en = dat_rsp_l2_pvld & _T_2124; // @[NV_NVDLA_CSC_dl_for_check.scala 1100:41:@1739.4]
  assign _GEN_149 = dat_rsp_sft_d1_en ? dat_rsp_l0_sft : {{256'd0}, dat_rsp_l0_sft_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:24:@1740.4]
  assign _GEN_150 = dat_rsp_sft_d2_en ? dat_rsp_l0_sft_d1 : {{128'd0}, dat_rsp_l0_sft_d2}; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1743.4]
  assign _GEN_151 = dat_rsp_sft_d2_en ? dat_rsp_l1_sft : {{384'd0}, dat_rsp_l1_sft_d2}; // @[NV_NVDLA_CSC_dl_for_check.scala 1105:24:@1743.4]
  assign _GEN_154 = dat_rsp_sft_d3_en ? dat_rsp_l2_sft : {{384'd0}, dat_rsp_l2_sft_d3}; // @[NV_NVDLA_CSC_dl_for_check.scala 1109:24:@1747.4]
  assign _T_2132 = 319'hffffffffffffffff << dat_rsp_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:56:@1753.4]
  assign _T_2133 = _T_2132[63:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:73:@1754.4]
  assign dat_rsp_ori_mask = ~ _T_2133; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:24:@1755.4]
  assign _T_2135 = dat_rsp_cur_sub_h >= 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:51:@1756.4]
  assign dat_rsp_cur_h_mask_p1 = _T_2135 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:32:@1758.4]
  assign _T_2143 = dat_rsp_cur_sub_h >= 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:51:@1759.4]
  assign dat_rsp_cur_h_mask_p2 = _T_2143 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:32:@1761.4]
  assign _T_2151 = dat_rsp_cur_sub_h == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:51:@1762.4]
  assign dat_rsp_cur_h_mask_p3 = _T_2151 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:32:@1764.4]
  assign _T_2158 = dat_rsp_cur_h_mask_p1[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1124:57:@1765.4]
  assign dat_rsp_cur_h_e2_mask_8b = {_T_2158,32'hffffffff}; // @[Cat.scala 30:58:@1767.4]
  assign _T_2164 = dat_rsp_cur_h_mask_p3[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:57:@1768.4]
  assign _T_2165 = dat_rsp_cur_h_mask_p2[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:106:@1769.4]
  assign _T_2166 = dat_rsp_cur_h_mask_p1[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:155:@1770.4]
  assign dat_rsp_cur_h_e4_mask_8b = {_T_2164,_T_2165,_T_2166,16'hffff}; // @[Cat.scala 30:58:@1774.4]
  assign _T_2175 = sub_h_total_g11 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:43:@1775.4]
  assign _T_2176 = dat_rsp_ori_mask[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:89:@1776.4]
  assign _T_2178 = {_T_2176,_T_2176,_T_2176,_T_2176}; // @[Cat.scala 30:58:@1778.4]
  assign _T_2179 = _T_2178 & dat_rsp_cur_h_e4_mask_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:116:@1779.4]
  assign _T_2181 = sub_h_total_g11 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:43:@1780.4]
  assign _T_2182 = dat_rsp_ori_mask[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:89:@1781.4]
  assign _T_2183 = {_T_2182,_T_2182}; // @[Cat.scala 30:58:@1782.4]
  assign _T_2184 = _T_2183 & dat_rsp_cur_h_e2_mask_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:116:@1783.4]
  assign _T_2185 = _T_2181 ? _T_2184 : dat_rsp_ori_mask; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:26:@1784.4]
  assign dat_rsp_mask_8b = _T_2175 ? _T_2179 : _T_2185; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:26:@1785.4]
  assign _T_2186 = is_img_d1[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:35:@1786.4]
  assign dat_rsp_data_w_0 = _T_2186 ? dat_rsp_img_0 : dat_rsp_conv_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_1 = _T_2186 ? dat_rsp_img_1 : dat_rsp_conv_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_2 = _T_2186 ? dat_rsp_img_2 : dat_rsp_conv_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_3 = _T_2186 ? dat_rsp_img_3 : dat_rsp_conv_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_4 = _T_2186 ? dat_rsp_img_4 : dat_rsp_conv_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_5 = _T_2186 ? dat_rsp_img_5 : dat_rsp_conv_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_6 = _T_2186 ? dat_rsp_img_6 : dat_rsp_conv_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_7 = _T_2186 ? dat_rsp_img_7 : dat_rsp_conv_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_8 = _T_2186 ? dat_rsp_img_8 : dat_rsp_conv_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_9 = _T_2186 ? dat_rsp_img_9 : dat_rsp_conv_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_10 = _T_2186 ? dat_rsp_img_10 : dat_rsp_conv_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_11 = _T_2186 ? dat_rsp_img_11 : dat_rsp_conv_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_12 = _T_2186 ? dat_rsp_img_12 : dat_rsp_conv_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_13 = _T_2186 ? dat_rsp_img_13 : dat_rsp_conv_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_14 = _T_2186 ? dat_rsp_img_14 : dat_rsp_conv_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_15 = _T_2186 ? dat_rsp_img_15 : dat_rsp_conv_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_16 = _T_2186 ? dat_rsp_img_16 : dat_rsp_conv_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_17 = _T_2186 ? dat_rsp_img_17 : dat_rsp_conv_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_18 = _T_2186 ? dat_rsp_img_18 : dat_rsp_conv_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_19 = _T_2186 ? dat_rsp_img_19 : dat_rsp_conv_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_20 = _T_2186 ? dat_rsp_img_20 : dat_rsp_conv_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_21 = _T_2186 ? dat_rsp_img_21 : dat_rsp_conv_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_22 = _T_2186 ? dat_rsp_img_22 : dat_rsp_conv_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_23 = _T_2186 ? dat_rsp_img_23 : dat_rsp_conv_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_24 = _T_2186 ? dat_rsp_img_24 : dat_rsp_conv_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_25 = _T_2186 ? dat_rsp_img_25 : dat_rsp_conv_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_26 = _T_2186 ? dat_rsp_img_26 : dat_rsp_conv_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_27 = _T_2186 ? dat_rsp_img_27 : dat_rsp_conv_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_28 = _T_2186 ? dat_rsp_img_28 : dat_rsp_conv_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_29 = _T_2186 ? dat_rsp_img_29 : dat_rsp_conv_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_30 = _T_2186 ? dat_rsp_img_30 : dat_rsp_conv_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_31 = _T_2186 ? dat_rsp_img_31 : dat_rsp_conv_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_32 = _T_2186 ? dat_rsp_img_32 : dat_rsp_conv_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_33 = _T_2186 ? dat_rsp_img_33 : dat_rsp_conv_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_34 = _T_2186 ? dat_rsp_img_34 : dat_rsp_conv_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_35 = _T_2186 ? dat_rsp_img_35 : dat_rsp_conv_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_36 = _T_2186 ? dat_rsp_img_36 : dat_rsp_conv_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_37 = _T_2186 ? dat_rsp_img_37 : dat_rsp_conv_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_38 = _T_2186 ? dat_rsp_img_38 : dat_rsp_conv_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_39 = _T_2186 ? dat_rsp_img_39 : dat_rsp_conv_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_40 = _T_2186 ? dat_rsp_img_40 : dat_rsp_conv_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_41 = _T_2186 ? dat_rsp_img_41 : dat_rsp_conv_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_42 = _T_2186 ? dat_rsp_img_42 : dat_rsp_conv_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_43 = _T_2186 ? dat_rsp_img_43 : dat_rsp_conv_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_44 = _T_2186 ? dat_rsp_img_44 : dat_rsp_conv_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_45 = _T_2186 ? dat_rsp_img_45 : dat_rsp_conv_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_46 = _T_2186 ? dat_rsp_img_46 : dat_rsp_conv_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_47 = _T_2186 ? dat_rsp_img_47 : dat_rsp_conv_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_48 = _T_2186 ? dat_rsp_img_48 : dat_rsp_conv_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_49 = _T_2186 ? dat_rsp_img_49 : dat_rsp_conv_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_50 = _T_2186 ? dat_rsp_img_50 : dat_rsp_conv_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_51 = _T_2186 ? dat_rsp_img_51 : dat_rsp_conv_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_52 = _T_2186 ? dat_rsp_img_52 : dat_rsp_conv_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_53 = _T_2186 ? dat_rsp_img_53 : dat_rsp_conv_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_54 = _T_2186 ? dat_rsp_img_54 : dat_rsp_conv_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_55 = _T_2186 ? dat_rsp_img_55 : dat_rsp_conv_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_56 = _T_2186 ? dat_rsp_img_56 : dat_rsp_conv_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_57 = _T_2186 ? dat_rsp_img_57 : dat_rsp_conv_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_58 = _T_2186 ? dat_rsp_img_58 : dat_rsp_conv_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_59 = _T_2186 ? dat_rsp_img_59 : dat_rsp_conv_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_60 = _T_2186 ? dat_rsp_img_60 : dat_rsp_conv_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_61 = _T_2186 ? dat_rsp_img_61 : dat_rsp_conv_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_62 = _T_2186 ? dat_rsp_img_62 : dat_rsp_conv_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_data_w_63 = _T_2186 ? dat_rsp_img_63 : dat_rsp_conv_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1132:25:@1787.4]
  assign dat_rsp_mask_val_int8_0 = dat_rsp_data_w_0 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1788.4]
  assign dat_rsp_mask_val_int8_1 = dat_rsp_data_w_1 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1789.4]
  assign dat_rsp_mask_val_int8_2 = dat_rsp_data_w_2 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1790.4]
  assign dat_rsp_mask_val_int8_3 = dat_rsp_data_w_3 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1791.4]
  assign dat_rsp_mask_val_int8_4 = dat_rsp_data_w_4 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1792.4]
  assign dat_rsp_mask_val_int8_5 = dat_rsp_data_w_5 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1793.4]
  assign dat_rsp_mask_val_int8_6 = dat_rsp_data_w_6 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1794.4]
  assign dat_rsp_mask_val_int8_7 = dat_rsp_data_w_7 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1795.4]
  assign dat_rsp_mask_val_int8_8 = dat_rsp_data_w_8 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1796.4]
  assign dat_rsp_mask_val_int8_9 = dat_rsp_data_w_9 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1797.4]
  assign dat_rsp_mask_val_int8_10 = dat_rsp_data_w_10 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1798.4]
  assign dat_rsp_mask_val_int8_11 = dat_rsp_data_w_11 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1799.4]
  assign dat_rsp_mask_val_int8_12 = dat_rsp_data_w_12 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1800.4]
  assign dat_rsp_mask_val_int8_13 = dat_rsp_data_w_13 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1801.4]
  assign dat_rsp_mask_val_int8_14 = dat_rsp_data_w_14 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1802.4]
  assign dat_rsp_mask_val_int8_15 = dat_rsp_data_w_15 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1803.4]
  assign dat_rsp_mask_val_int8_16 = dat_rsp_data_w_16 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1804.4]
  assign dat_rsp_mask_val_int8_17 = dat_rsp_data_w_17 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1805.4]
  assign dat_rsp_mask_val_int8_18 = dat_rsp_data_w_18 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1806.4]
  assign dat_rsp_mask_val_int8_19 = dat_rsp_data_w_19 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1807.4]
  assign dat_rsp_mask_val_int8_20 = dat_rsp_data_w_20 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1808.4]
  assign dat_rsp_mask_val_int8_21 = dat_rsp_data_w_21 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1809.4]
  assign dat_rsp_mask_val_int8_22 = dat_rsp_data_w_22 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1810.4]
  assign dat_rsp_mask_val_int8_23 = dat_rsp_data_w_23 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1811.4]
  assign dat_rsp_mask_val_int8_24 = dat_rsp_data_w_24 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1812.4]
  assign dat_rsp_mask_val_int8_25 = dat_rsp_data_w_25 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1813.4]
  assign dat_rsp_mask_val_int8_26 = dat_rsp_data_w_26 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1814.4]
  assign dat_rsp_mask_val_int8_27 = dat_rsp_data_w_27 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1815.4]
  assign dat_rsp_mask_val_int8_28 = dat_rsp_data_w_28 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1816.4]
  assign dat_rsp_mask_val_int8_29 = dat_rsp_data_w_29 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1817.4]
  assign dat_rsp_mask_val_int8_30 = dat_rsp_data_w_30 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1818.4]
  assign dat_rsp_mask_val_int8_31 = dat_rsp_data_w_31 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1819.4]
  assign dat_rsp_mask_val_int8_32 = dat_rsp_data_w_32 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1820.4]
  assign dat_rsp_mask_val_int8_33 = dat_rsp_data_w_33 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1821.4]
  assign dat_rsp_mask_val_int8_34 = dat_rsp_data_w_34 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1822.4]
  assign dat_rsp_mask_val_int8_35 = dat_rsp_data_w_35 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1823.4]
  assign dat_rsp_mask_val_int8_36 = dat_rsp_data_w_36 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1824.4]
  assign dat_rsp_mask_val_int8_37 = dat_rsp_data_w_37 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1825.4]
  assign dat_rsp_mask_val_int8_38 = dat_rsp_data_w_38 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1826.4]
  assign dat_rsp_mask_val_int8_39 = dat_rsp_data_w_39 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1827.4]
  assign dat_rsp_mask_val_int8_40 = dat_rsp_data_w_40 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1828.4]
  assign dat_rsp_mask_val_int8_41 = dat_rsp_data_w_41 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1829.4]
  assign dat_rsp_mask_val_int8_42 = dat_rsp_data_w_42 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1830.4]
  assign dat_rsp_mask_val_int8_43 = dat_rsp_data_w_43 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1831.4]
  assign dat_rsp_mask_val_int8_44 = dat_rsp_data_w_44 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1832.4]
  assign dat_rsp_mask_val_int8_45 = dat_rsp_data_w_45 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1833.4]
  assign dat_rsp_mask_val_int8_46 = dat_rsp_data_w_46 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1834.4]
  assign dat_rsp_mask_val_int8_47 = dat_rsp_data_w_47 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1835.4]
  assign dat_rsp_mask_val_int8_48 = dat_rsp_data_w_48 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1836.4]
  assign dat_rsp_mask_val_int8_49 = dat_rsp_data_w_49 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1837.4]
  assign dat_rsp_mask_val_int8_50 = dat_rsp_data_w_50 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1838.4]
  assign dat_rsp_mask_val_int8_51 = dat_rsp_data_w_51 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1839.4]
  assign dat_rsp_mask_val_int8_52 = dat_rsp_data_w_52 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1840.4]
  assign dat_rsp_mask_val_int8_53 = dat_rsp_data_w_53 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1841.4]
  assign dat_rsp_mask_val_int8_54 = dat_rsp_data_w_54 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1842.4]
  assign dat_rsp_mask_val_int8_55 = dat_rsp_data_w_55 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1843.4]
  assign dat_rsp_mask_val_int8_56 = dat_rsp_data_w_56 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1844.4]
  assign dat_rsp_mask_val_int8_57 = dat_rsp_data_w_57 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1845.4]
  assign dat_rsp_mask_val_int8_58 = dat_rsp_data_w_58 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1846.4]
  assign dat_rsp_mask_val_int8_59 = dat_rsp_data_w_59 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1847.4]
  assign dat_rsp_mask_val_int8_60 = dat_rsp_data_w_60 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1848.4]
  assign dat_rsp_mask_val_int8_61 = dat_rsp_data_w_61 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1849.4]
  assign dat_rsp_mask_val_int8_62 = dat_rsp_data_w_62 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1850.4]
  assign dat_rsp_mask_val_int8_63 = dat_rsp_data_w_63 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:97:@1851.4]
  assign _T_2515 = dat_rsp_mask_8b[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1917.4]
  assign dat_rsp_mask_w_0 = _T_2515 & dat_rsp_mask_val_int8_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1918.4]
  assign _T_2517 = dat_rsp_mask_8b[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1919.4]
  assign dat_rsp_mask_w_1 = _T_2517 & dat_rsp_mask_val_int8_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1920.4]
  assign _T_2519 = dat_rsp_mask_8b[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1921.4]
  assign dat_rsp_mask_w_2 = _T_2519 & dat_rsp_mask_val_int8_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1922.4]
  assign _T_2521 = dat_rsp_mask_8b[3]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1923.4]
  assign dat_rsp_mask_w_3 = _T_2521 & dat_rsp_mask_val_int8_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1924.4]
  assign _T_2523 = dat_rsp_mask_8b[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1925.4]
  assign dat_rsp_mask_w_4 = _T_2523 & dat_rsp_mask_val_int8_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1926.4]
  assign _T_2525 = dat_rsp_mask_8b[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1927.4]
  assign dat_rsp_mask_w_5 = _T_2525 & dat_rsp_mask_val_int8_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1928.4]
  assign _T_2527 = dat_rsp_mask_8b[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1929.4]
  assign dat_rsp_mask_w_6 = _T_2527 & dat_rsp_mask_val_int8_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1930.4]
  assign _T_2529 = dat_rsp_mask_8b[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1931.4]
  assign dat_rsp_mask_w_7 = _T_2529 & dat_rsp_mask_val_int8_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1932.4]
  assign _T_2531 = dat_rsp_mask_8b[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1933.4]
  assign dat_rsp_mask_w_8 = _T_2531 & dat_rsp_mask_val_int8_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1934.4]
  assign _T_2533 = dat_rsp_mask_8b[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1935.4]
  assign dat_rsp_mask_w_9 = _T_2533 & dat_rsp_mask_val_int8_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1936.4]
  assign _T_2535 = dat_rsp_mask_8b[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1937.4]
  assign dat_rsp_mask_w_10 = _T_2535 & dat_rsp_mask_val_int8_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1938.4]
  assign _T_2537 = dat_rsp_mask_8b[11]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1939.4]
  assign dat_rsp_mask_w_11 = _T_2537 & dat_rsp_mask_val_int8_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1940.4]
  assign _T_2539 = dat_rsp_mask_8b[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1941.4]
  assign dat_rsp_mask_w_12 = _T_2539 & dat_rsp_mask_val_int8_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1942.4]
  assign _T_2541 = dat_rsp_mask_8b[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1943.4]
  assign dat_rsp_mask_w_13 = _T_2541 & dat_rsp_mask_val_int8_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1944.4]
  assign _T_2543 = dat_rsp_mask_8b[14]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1945.4]
  assign dat_rsp_mask_w_14 = _T_2543 & dat_rsp_mask_val_int8_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1946.4]
  assign _T_2545 = dat_rsp_mask_8b[15]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1947.4]
  assign dat_rsp_mask_w_15 = _T_2545 & dat_rsp_mask_val_int8_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1948.4]
  assign _T_2547 = dat_rsp_mask_8b[16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1949.4]
  assign dat_rsp_mask_w_16 = _T_2547 & dat_rsp_mask_val_int8_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1950.4]
  assign _T_2549 = dat_rsp_mask_8b[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1951.4]
  assign dat_rsp_mask_w_17 = _T_2549 & dat_rsp_mask_val_int8_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1952.4]
  assign _T_2551 = dat_rsp_mask_8b[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1953.4]
  assign dat_rsp_mask_w_18 = _T_2551 & dat_rsp_mask_val_int8_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1954.4]
  assign _T_2553 = dat_rsp_mask_8b[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1955.4]
  assign dat_rsp_mask_w_19 = _T_2553 & dat_rsp_mask_val_int8_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1956.4]
  assign _T_2555 = dat_rsp_mask_8b[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1957.4]
  assign dat_rsp_mask_w_20 = _T_2555 & dat_rsp_mask_val_int8_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1958.4]
  assign _T_2557 = dat_rsp_mask_8b[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1959.4]
  assign dat_rsp_mask_w_21 = _T_2557 & dat_rsp_mask_val_int8_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1960.4]
  assign _T_2559 = dat_rsp_mask_8b[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1961.4]
  assign dat_rsp_mask_w_22 = _T_2559 & dat_rsp_mask_val_int8_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1962.4]
  assign _T_2561 = dat_rsp_mask_8b[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1963.4]
  assign dat_rsp_mask_w_23 = _T_2561 & dat_rsp_mask_val_int8_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1964.4]
  assign _T_2563 = dat_rsp_mask_8b[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1965.4]
  assign dat_rsp_mask_w_24 = _T_2563 & dat_rsp_mask_val_int8_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1966.4]
  assign _T_2565 = dat_rsp_mask_8b[25]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1967.4]
  assign dat_rsp_mask_w_25 = _T_2565 & dat_rsp_mask_val_int8_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1968.4]
  assign _T_2567 = dat_rsp_mask_8b[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1969.4]
  assign dat_rsp_mask_w_26 = _T_2567 & dat_rsp_mask_val_int8_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1970.4]
  assign _T_2569 = dat_rsp_mask_8b[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1971.4]
  assign dat_rsp_mask_w_27 = _T_2569 & dat_rsp_mask_val_int8_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1972.4]
  assign _T_2571 = dat_rsp_mask_8b[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1973.4]
  assign dat_rsp_mask_w_28 = _T_2571 & dat_rsp_mask_val_int8_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1974.4]
  assign _T_2573 = dat_rsp_mask_8b[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1975.4]
  assign dat_rsp_mask_w_29 = _T_2573 & dat_rsp_mask_val_int8_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1976.4]
  assign _T_2575 = dat_rsp_mask_8b[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1977.4]
  assign dat_rsp_mask_w_30 = _T_2575 & dat_rsp_mask_val_int8_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1978.4]
  assign _T_2577 = dat_rsp_mask_8b[31]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1979.4]
  assign dat_rsp_mask_w_31 = _T_2577 & dat_rsp_mask_val_int8_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1980.4]
  assign _T_2579 = dat_rsp_mask_8b[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1981.4]
  assign dat_rsp_mask_w_32 = _T_2579 & dat_rsp_mask_val_int8_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1982.4]
  assign _T_2581 = dat_rsp_mask_8b[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1983.4]
  assign dat_rsp_mask_w_33 = _T_2581 & dat_rsp_mask_val_int8_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1984.4]
  assign _T_2583 = dat_rsp_mask_8b[34]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1985.4]
  assign dat_rsp_mask_w_34 = _T_2583 & dat_rsp_mask_val_int8_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1986.4]
  assign _T_2585 = dat_rsp_mask_8b[35]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1987.4]
  assign dat_rsp_mask_w_35 = _T_2585 & dat_rsp_mask_val_int8_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1988.4]
  assign _T_2587 = dat_rsp_mask_8b[36]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1989.4]
  assign dat_rsp_mask_w_36 = _T_2587 & dat_rsp_mask_val_int8_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1990.4]
  assign _T_2589 = dat_rsp_mask_8b[37]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1991.4]
  assign dat_rsp_mask_w_37 = _T_2589 & dat_rsp_mask_val_int8_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1992.4]
  assign _T_2591 = dat_rsp_mask_8b[38]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1993.4]
  assign dat_rsp_mask_w_38 = _T_2591 & dat_rsp_mask_val_int8_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1994.4]
  assign _T_2593 = dat_rsp_mask_8b[39]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1995.4]
  assign dat_rsp_mask_w_39 = _T_2593 & dat_rsp_mask_val_int8_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1996.4]
  assign _T_2595 = dat_rsp_mask_8b[40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1997.4]
  assign dat_rsp_mask_w_40 = _T_2595 & dat_rsp_mask_val_int8_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@1998.4]
  assign _T_2597 = dat_rsp_mask_8b[41]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@1999.4]
  assign dat_rsp_mask_w_41 = _T_2597 & dat_rsp_mask_val_int8_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2000.4]
  assign _T_2599 = dat_rsp_mask_8b[42]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2001.4]
  assign dat_rsp_mask_w_42 = _T_2599 & dat_rsp_mask_val_int8_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2002.4]
  assign _T_2601 = dat_rsp_mask_8b[43]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2003.4]
  assign dat_rsp_mask_w_43 = _T_2601 & dat_rsp_mask_val_int8_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2004.4]
  assign _T_2603 = dat_rsp_mask_8b[44]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2005.4]
  assign dat_rsp_mask_w_44 = _T_2603 & dat_rsp_mask_val_int8_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2006.4]
  assign _T_2605 = dat_rsp_mask_8b[45]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2007.4]
  assign dat_rsp_mask_w_45 = _T_2605 & dat_rsp_mask_val_int8_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2008.4]
  assign _T_2607 = dat_rsp_mask_8b[46]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2009.4]
  assign dat_rsp_mask_w_46 = _T_2607 & dat_rsp_mask_val_int8_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2010.4]
  assign _T_2609 = dat_rsp_mask_8b[47]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2011.4]
  assign dat_rsp_mask_w_47 = _T_2609 & dat_rsp_mask_val_int8_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2012.4]
  assign _T_2611 = dat_rsp_mask_8b[48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2013.4]
  assign dat_rsp_mask_w_48 = _T_2611 & dat_rsp_mask_val_int8_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2014.4]
  assign _T_2613 = dat_rsp_mask_8b[49]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2015.4]
  assign dat_rsp_mask_w_49 = _T_2613 & dat_rsp_mask_val_int8_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2016.4]
  assign _T_2615 = dat_rsp_mask_8b[50]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2017.4]
  assign dat_rsp_mask_w_50 = _T_2615 & dat_rsp_mask_val_int8_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2018.4]
  assign _T_2617 = dat_rsp_mask_8b[51]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2019.4]
  assign dat_rsp_mask_w_51 = _T_2617 & dat_rsp_mask_val_int8_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2020.4]
  assign _T_2619 = dat_rsp_mask_8b[52]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2021.4]
  assign dat_rsp_mask_w_52 = _T_2619 & dat_rsp_mask_val_int8_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2022.4]
  assign _T_2621 = dat_rsp_mask_8b[53]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2023.4]
  assign dat_rsp_mask_w_53 = _T_2621 & dat_rsp_mask_val_int8_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2024.4]
  assign _T_2623 = dat_rsp_mask_8b[54]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2025.4]
  assign dat_rsp_mask_w_54 = _T_2623 & dat_rsp_mask_val_int8_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2026.4]
  assign _T_2625 = dat_rsp_mask_8b[55]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2027.4]
  assign dat_rsp_mask_w_55 = _T_2625 & dat_rsp_mask_val_int8_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2028.4]
  assign _T_2627 = dat_rsp_mask_8b[56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2029.4]
  assign dat_rsp_mask_w_56 = _T_2627 & dat_rsp_mask_val_int8_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2030.4]
  assign _T_2629 = dat_rsp_mask_8b[57]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2031.4]
  assign dat_rsp_mask_w_57 = _T_2629 & dat_rsp_mask_val_int8_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2032.4]
  assign _T_2631 = dat_rsp_mask_8b[58]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2033.4]
  assign dat_rsp_mask_w_58 = _T_2631 & dat_rsp_mask_val_int8_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2034.4]
  assign _T_2633 = dat_rsp_mask_8b[59]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2035.4]
  assign dat_rsp_mask_w_59 = _T_2633 & dat_rsp_mask_val_int8_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2036.4]
  assign _T_2635 = dat_rsp_mask_8b[60]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2037.4]
  assign dat_rsp_mask_w_60 = _T_2635 & dat_rsp_mask_val_int8_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2038.4]
  assign _T_2637 = dat_rsp_mask_8b[61]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2039.4]
  assign dat_rsp_mask_w_61 = _T_2637 & dat_rsp_mask_val_int8_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2040.4]
  assign _T_2639 = dat_rsp_mask_8b[62]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2041.4]
  assign dat_rsp_mask_w_62 = _T_2639 & dat_rsp_mask_val_int8_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2042.4]
  assign _T_2641 = dat_rsp_mask_8b[63]; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:80:@2043.4]
  assign dat_rsp_mask_w_63 = _T_2641 & dat_rsp_mask_val_int8_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:83:@2044.4]
  assign _GEN_155 = dat_rsp_pvld ? dat_rsp_flag : dat_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1154:21:@2180.4]
  assign _GEN_156 = dat_rsp_pvld ? dat_rsp_mask_w_0 : dat_out_bypass_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_157 = dat_rsp_pvld ? dat_rsp_mask_w_1 : dat_out_bypass_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_158 = dat_rsp_pvld ? dat_rsp_mask_w_2 : dat_out_bypass_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_159 = dat_rsp_pvld ? dat_rsp_mask_w_3 : dat_out_bypass_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_160 = dat_rsp_pvld ? dat_rsp_mask_w_4 : dat_out_bypass_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_161 = dat_rsp_pvld ? dat_rsp_mask_w_5 : dat_out_bypass_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_162 = dat_rsp_pvld ? dat_rsp_mask_w_6 : dat_out_bypass_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_163 = dat_rsp_pvld ? dat_rsp_mask_w_7 : dat_out_bypass_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_164 = dat_rsp_pvld ? dat_rsp_mask_w_8 : dat_out_bypass_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_165 = dat_rsp_pvld ? dat_rsp_mask_w_9 : dat_out_bypass_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_166 = dat_rsp_pvld ? dat_rsp_mask_w_10 : dat_out_bypass_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_167 = dat_rsp_pvld ? dat_rsp_mask_w_11 : dat_out_bypass_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_168 = dat_rsp_pvld ? dat_rsp_mask_w_12 : dat_out_bypass_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_169 = dat_rsp_pvld ? dat_rsp_mask_w_13 : dat_out_bypass_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_170 = dat_rsp_pvld ? dat_rsp_mask_w_14 : dat_out_bypass_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_171 = dat_rsp_pvld ? dat_rsp_mask_w_15 : dat_out_bypass_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_172 = dat_rsp_pvld ? dat_rsp_mask_w_16 : dat_out_bypass_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_173 = dat_rsp_pvld ? dat_rsp_mask_w_17 : dat_out_bypass_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_174 = dat_rsp_pvld ? dat_rsp_mask_w_18 : dat_out_bypass_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_175 = dat_rsp_pvld ? dat_rsp_mask_w_19 : dat_out_bypass_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_176 = dat_rsp_pvld ? dat_rsp_mask_w_20 : dat_out_bypass_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_177 = dat_rsp_pvld ? dat_rsp_mask_w_21 : dat_out_bypass_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_178 = dat_rsp_pvld ? dat_rsp_mask_w_22 : dat_out_bypass_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_179 = dat_rsp_pvld ? dat_rsp_mask_w_23 : dat_out_bypass_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_180 = dat_rsp_pvld ? dat_rsp_mask_w_24 : dat_out_bypass_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_181 = dat_rsp_pvld ? dat_rsp_mask_w_25 : dat_out_bypass_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_182 = dat_rsp_pvld ? dat_rsp_mask_w_26 : dat_out_bypass_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_183 = dat_rsp_pvld ? dat_rsp_mask_w_27 : dat_out_bypass_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_184 = dat_rsp_pvld ? dat_rsp_mask_w_28 : dat_out_bypass_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_185 = dat_rsp_pvld ? dat_rsp_mask_w_29 : dat_out_bypass_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_186 = dat_rsp_pvld ? dat_rsp_mask_w_30 : dat_out_bypass_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_187 = dat_rsp_pvld ? dat_rsp_mask_w_31 : dat_out_bypass_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_188 = dat_rsp_pvld ? dat_rsp_mask_w_32 : dat_out_bypass_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_189 = dat_rsp_pvld ? dat_rsp_mask_w_33 : dat_out_bypass_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_190 = dat_rsp_pvld ? dat_rsp_mask_w_34 : dat_out_bypass_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_191 = dat_rsp_pvld ? dat_rsp_mask_w_35 : dat_out_bypass_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_192 = dat_rsp_pvld ? dat_rsp_mask_w_36 : dat_out_bypass_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_193 = dat_rsp_pvld ? dat_rsp_mask_w_37 : dat_out_bypass_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_194 = dat_rsp_pvld ? dat_rsp_mask_w_38 : dat_out_bypass_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_195 = dat_rsp_pvld ? dat_rsp_mask_w_39 : dat_out_bypass_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_196 = dat_rsp_pvld ? dat_rsp_mask_w_40 : dat_out_bypass_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_197 = dat_rsp_pvld ? dat_rsp_mask_w_41 : dat_out_bypass_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_198 = dat_rsp_pvld ? dat_rsp_mask_w_42 : dat_out_bypass_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_199 = dat_rsp_pvld ? dat_rsp_mask_w_43 : dat_out_bypass_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_200 = dat_rsp_pvld ? dat_rsp_mask_w_44 : dat_out_bypass_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_201 = dat_rsp_pvld ? dat_rsp_mask_w_45 : dat_out_bypass_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_202 = dat_rsp_pvld ? dat_rsp_mask_w_46 : dat_out_bypass_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_203 = dat_rsp_pvld ? dat_rsp_mask_w_47 : dat_out_bypass_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_204 = dat_rsp_pvld ? dat_rsp_mask_w_48 : dat_out_bypass_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_205 = dat_rsp_pvld ? dat_rsp_mask_w_49 : dat_out_bypass_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_206 = dat_rsp_pvld ? dat_rsp_mask_w_50 : dat_out_bypass_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_207 = dat_rsp_pvld ? dat_rsp_mask_w_51 : dat_out_bypass_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_208 = dat_rsp_pvld ? dat_rsp_mask_w_52 : dat_out_bypass_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_209 = dat_rsp_pvld ? dat_rsp_mask_w_53 : dat_out_bypass_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_210 = dat_rsp_pvld ? dat_rsp_mask_w_54 : dat_out_bypass_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_211 = dat_rsp_pvld ? dat_rsp_mask_w_55 : dat_out_bypass_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_212 = dat_rsp_pvld ? dat_rsp_mask_w_56 : dat_out_bypass_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_213 = dat_rsp_pvld ? dat_rsp_mask_w_57 : dat_out_bypass_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_214 = dat_rsp_pvld ? dat_rsp_mask_w_58 : dat_out_bypass_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_215 = dat_rsp_pvld ? dat_rsp_mask_w_59 : dat_out_bypass_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_216 = dat_rsp_pvld ? dat_rsp_mask_w_60 : dat_out_bypass_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_217 = dat_rsp_pvld ? dat_rsp_mask_w_61 : dat_out_bypass_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_218 = dat_rsp_pvld ? dat_rsp_mask_w_62 : dat_out_bypass_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _GEN_219 = dat_rsp_pvld ? dat_rsp_mask_w_63 : dat_out_bypass_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1157:30:@2183.4]
  assign _T_3247 = dat_rsp_pvld & dat_rsp_mask_w_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2249.4]
  assign _T_3248 = dat_rsp_pvld & dat_rsp_mask_w_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2253.4]
  assign _T_3249 = dat_rsp_pvld & dat_rsp_mask_w_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2257.4]
  assign _T_3250 = dat_rsp_pvld & dat_rsp_mask_w_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2261.4]
  assign _T_3251 = dat_rsp_pvld & dat_rsp_mask_w_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2265.4]
  assign _T_3252 = dat_rsp_pvld & dat_rsp_mask_w_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2269.4]
  assign _T_3253 = dat_rsp_pvld & dat_rsp_mask_w_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2273.4]
  assign _T_3254 = dat_rsp_pvld & dat_rsp_mask_w_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2277.4]
  assign _T_3255 = dat_rsp_pvld & dat_rsp_mask_w_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2281.4]
  assign _T_3256 = dat_rsp_pvld & dat_rsp_mask_w_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2285.4]
  assign _T_3257 = dat_rsp_pvld & dat_rsp_mask_w_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2289.4]
  assign _T_3258 = dat_rsp_pvld & dat_rsp_mask_w_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2293.4]
  assign _T_3259 = dat_rsp_pvld & dat_rsp_mask_w_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2297.4]
  assign _T_3260 = dat_rsp_pvld & dat_rsp_mask_w_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2301.4]
  assign _T_3261 = dat_rsp_pvld & dat_rsp_mask_w_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2305.4]
  assign _T_3262 = dat_rsp_pvld & dat_rsp_mask_w_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2309.4]
  assign _T_3263 = dat_rsp_pvld & dat_rsp_mask_w_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2313.4]
  assign _T_3264 = dat_rsp_pvld & dat_rsp_mask_w_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2317.4]
  assign _T_3265 = dat_rsp_pvld & dat_rsp_mask_w_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2321.4]
  assign _T_3266 = dat_rsp_pvld & dat_rsp_mask_w_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2325.4]
  assign _T_3267 = dat_rsp_pvld & dat_rsp_mask_w_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2329.4]
  assign _T_3268 = dat_rsp_pvld & dat_rsp_mask_w_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2333.4]
  assign _T_3269 = dat_rsp_pvld & dat_rsp_mask_w_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2337.4]
  assign _T_3270 = dat_rsp_pvld & dat_rsp_mask_w_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2341.4]
  assign _T_3271 = dat_rsp_pvld & dat_rsp_mask_w_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2345.4]
  assign _T_3272 = dat_rsp_pvld & dat_rsp_mask_w_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2349.4]
  assign _T_3273 = dat_rsp_pvld & dat_rsp_mask_w_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2353.4]
  assign _T_3274 = dat_rsp_pvld & dat_rsp_mask_w_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2357.4]
  assign _T_3275 = dat_rsp_pvld & dat_rsp_mask_w_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2361.4]
  assign _T_3276 = dat_rsp_pvld & dat_rsp_mask_w_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2365.4]
  assign _T_3277 = dat_rsp_pvld & dat_rsp_mask_w_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2369.4]
  assign _T_3278 = dat_rsp_pvld & dat_rsp_mask_w_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2373.4]
  assign _T_3279 = dat_rsp_pvld & dat_rsp_mask_w_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2377.4]
  assign _T_3280 = dat_rsp_pvld & dat_rsp_mask_w_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2381.4]
  assign _T_3281 = dat_rsp_pvld & dat_rsp_mask_w_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2385.4]
  assign _T_3282 = dat_rsp_pvld & dat_rsp_mask_w_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2389.4]
  assign _T_3283 = dat_rsp_pvld & dat_rsp_mask_w_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2393.4]
  assign _T_3284 = dat_rsp_pvld & dat_rsp_mask_w_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2397.4]
  assign _T_3285 = dat_rsp_pvld & dat_rsp_mask_w_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2401.4]
  assign _T_3286 = dat_rsp_pvld & dat_rsp_mask_w_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2405.4]
  assign _T_3287 = dat_rsp_pvld & dat_rsp_mask_w_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2409.4]
  assign _T_3288 = dat_rsp_pvld & dat_rsp_mask_w_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2413.4]
  assign _T_3289 = dat_rsp_pvld & dat_rsp_mask_w_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2417.4]
  assign _T_3290 = dat_rsp_pvld & dat_rsp_mask_w_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2421.4]
  assign _T_3291 = dat_rsp_pvld & dat_rsp_mask_w_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2425.4]
  assign _T_3292 = dat_rsp_pvld & dat_rsp_mask_w_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2429.4]
  assign _T_3293 = dat_rsp_pvld & dat_rsp_mask_w_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2433.4]
  assign _T_3294 = dat_rsp_pvld & dat_rsp_mask_w_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2437.4]
  assign _T_3295 = dat_rsp_pvld & dat_rsp_mask_w_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2441.4]
  assign _T_3296 = dat_rsp_pvld & dat_rsp_mask_w_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2445.4]
  assign _T_3297 = dat_rsp_pvld & dat_rsp_mask_w_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2449.4]
  assign _T_3298 = dat_rsp_pvld & dat_rsp_mask_w_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2453.4]
  assign _T_3299 = dat_rsp_pvld & dat_rsp_mask_w_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2457.4]
  assign _T_3300 = dat_rsp_pvld & dat_rsp_mask_w_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2461.4]
  assign _T_3301 = dat_rsp_pvld & dat_rsp_mask_w_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2465.4]
  assign _T_3302 = dat_rsp_pvld & dat_rsp_mask_w_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2469.4]
  assign _T_3303 = dat_rsp_pvld & dat_rsp_mask_w_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2473.4]
  assign _T_3304 = dat_rsp_pvld & dat_rsp_mask_w_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2477.4]
  assign _T_3305 = dat_rsp_pvld & dat_rsp_mask_w_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2481.4]
  assign _T_3306 = dat_rsp_pvld & dat_rsp_mask_w_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2485.4]
  assign _T_3307 = dat_rsp_pvld & dat_rsp_mask_w_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2489.4]
  assign _T_3308 = dat_rsp_pvld & dat_rsp_mask_w_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2493.4]
  assign _T_3309 = dat_rsp_pvld & dat_rsp_mask_w_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2497.4]
  assign _T_3310 = dat_rsp_pvld & dat_rsp_mask_w_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:34:@2501.4]
  assign _T_3846 = ~ dat_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:24:@2574.4]
  assign dat_out_mask_0 = _T_3846 ? 1'h0 : dat_out_bypass_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_1 = _T_3846 ? 1'h0 : dat_out_bypass_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_2 = _T_3846 ? 1'h0 : dat_out_bypass_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_3 = _T_3846 ? 1'h0 : dat_out_bypass_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_4 = _T_3846 ? 1'h0 : dat_out_bypass_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_5 = _T_3846 ? 1'h0 : dat_out_bypass_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_6 = _T_3846 ? 1'h0 : dat_out_bypass_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_7 = _T_3846 ? 1'h0 : dat_out_bypass_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_8 = _T_3846 ? 1'h0 : dat_out_bypass_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_9 = _T_3846 ? 1'h0 : dat_out_bypass_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_10 = _T_3846 ? 1'h0 : dat_out_bypass_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_11 = _T_3846 ? 1'h0 : dat_out_bypass_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_12 = _T_3846 ? 1'h0 : dat_out_bypass_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_13 = _T_3846 ? 1'h0 : dat_out_bypass_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_14 = _T_3846 ? 1'h0 : dat_out_bypass_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_15 = _T_3846 ? 1'h0 : dat_out_bypass_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_16 = _T_3846 ? 1'h0 : dat_out_bypass_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_17 = _T_3846 ? 1'h0 : dat_out_bypass_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_18 = _T_3846 ? 1'h0 : dat_out_bypass_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_19 = _T_3846 ? 1'h0 : dat_out_bypass_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_20 = _T_3846 ? 1'h0 : dat_out_bypass_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_21 = _T_3846 ? 1'h0 : dat_out_bypass_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_22 = _T_3846 ? 1'h0 : dat_out_bypass_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_23 = _T_3846 ? 1'h0 : dat_out_bypass_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_24 = _T_3846 ? 1'h0 : dat_out_bypass_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_25 = _T_3846 ? 1'h0 : dat_out_bypass_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_26 = _T_3846 ? 1'h0 : dat_out_bypass_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_27 = _T_3846 ? 1'h0 : dat_out_bypass_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_28 = _T_3846 ? 1'h0 : dat_out_bypass_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_29 = _T_3846 ? 1'h0 : dat_out_bypass_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_30 = _T_3846 ? 1'h0 : dat_out_bypass_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_31 = _T_3846 ? 1'h0 : dat_out_bypass_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_32 = _T_3846 ? 1'h0 : dat_out_bypass_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_33 = _T_3846 ? 1'h0 : dat_out_bypass_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_34 = _T_3846 ? 1'h0 : dat_out_bypass_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_35 = _T_3846 ? 1'h0 : dat_out_bypass_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_36 = _T_3846 ? 1'h0 : dat_out_bypass_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_37 = _T_3846 ? 1'h0 : dat_out_bypass_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_38 = _T_3846 ? 1'h0 : dat_out_bypass_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_39 = _T_3846 ? 1'h0 : dat_out_bypass_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_40 = _T_3846 ? 1'h0 : dat_out_bypass_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_41 = _T_3846 ? 1'h0 : dat_out_bypass_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_42 = _T_3846 ? 1'h0 : dat_out_bypass_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_43 = _T_3846 ? 1'h0 : dat_out_bypass_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_44 = _T_3846 ? 1'h0 : dat_out_bypass_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_45 = _T_3846 ? 1'h0 : dat_out_bypass_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_46 = _T_3846 ? 1'h0 : dat_out_bypass_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_47 = _T_3846 ? 1'h0 : dat_out_bypass_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_48 = _T_3846 ? 1'h0 : dat_out_bypass_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_49 = _T_3846 ? 1'h0 : dat_out_bypass_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_50 = _T_3846 ? 1'h0 : dat_out_bypass_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_51 = _T_3846 ? 1'h0 : dat_out_bypass_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_52 = _T_3846 ? 1'h0 : dat_out_bypass_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_53 = _T_3846 ? 1'h0 : dat_out_bypass_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_54 = _T_3846 ? 1'h0 : dat_out_bypass_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_55 = _T_3846 ? 1'h0 : dat_out_bypass_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_56 = _T_3846 ? 1'h0 : dat_out_bypass_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_57 = _T_3846 ? 1'h0 : dat_out_bypass_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_58 = _T_3846 ? 1'h0 : dat_out_bypass_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_59 = _T_3846 ? 1'h0 : dat_out_bypass_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_60 = _T_3846 ? 1'h0 : dat_out_bypass_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_61 = _T_3846 ? 1'h0 : dat_out_bypass_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_62 = _T_3846 ? 1'h0 : dat_out_bypass_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign dat_out_mask_63 = _T_3846 ? 1'h0 : dat_out_bypass_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1175:23:@2640.4]
  assign _T_4112 = dat_out_pvld | dl_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:19:@2642.4]
  assign _GEN_284 = _T_4112 ? dat_out_mask_0 : dl_out_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_285 = _T_4112 ? dat_out_mask_1 : dl_out_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_286 = _T_4112 ? dat_out_mask_2 : dl_out_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_287 = _T_4112 ? dat_out_mask_3 : dl_out_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_288 = _T_4112 ? dat_out_mask_4 : dl_out_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_289 = _T_4112 ? dat_out_mask_5 : dl_out_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_290 = _T_4112 ? dat_out_mask_6 : dl_out_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_291 = _T_4112 ? dat_out_mask_7 : dl_out_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_292 = _T_4112 ? dat_out_mask_8 : dl_out_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_293 = _T_4112 ? dat_out_mask_9 : dl_out_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_294 = _T_4112 ? dat_out_mask_10 : dl_out_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_295 = _T_4112 ? dat_out_mask_11 : dl_out_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_296 = _T_4112 ? dat_out_mask_12 : dl_out_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_297 = _T_4112 ? dat_out_mask_13 : dl_out_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_298 = _T_4112 ? dat_out_mask_14 : dl_out_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_299 = _T_4112 ? dat_out_mask_15 : dl_out_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_300 = _T_4112 ? dat_out_mask_16 : dl_out_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_301 = _T_4112 ? dat_out_mask_17 : dl_out_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_302 = _T_4112 ? dat_out_mask_18 : dl_out_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_303 = _T_4112 ? dat_out_mask_19 : dl_out_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_304 = _T_4112 ? dat_out_mask_20 : dl_out_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_305 = _T_4112 ? dat_out_mask_21 : dl_out_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_306 = _T_4112 ? dat_out_mask_22 : dl_out_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_307 = _T_4112 ? dat_out_mask_23 : dl_out_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_308 = _T_4112 ? dat_out_mask_24 : dl_out_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_309 = _T_4112 ? dat_out_mask_25 : dl_out_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_310 = _T_4112 ? dat_out_mask_26 : dl_out_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_311 = _T_4112 ? dat_out_mask_27 : dl_out_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_312 = _T_4112 ? dat_out_mask_28 : dl_out_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_313 = _T_4112 ? dat_out_mask_29 : dl_out_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_314 = _T_4112 ? dat_out_mask_30 : dl_out_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_315 = _T_4112 ? dat_out_mask_31 : dl_out_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_316 = _T_4112 ? dat_out_mask_32 : dl_out_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_317 = _T_4112 ? dat_out_mask_33 : dl_out_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_318 = _T_4112 ? dat_out_mask_34 : dl_out_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_319 = _T_4112 ? dat_out_mask_35 : dl_out_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_320 = _T_4112 ? dat_out_mask_36 : dl_out_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_321 = _T_4112 ? dat_out_mask_37 : dl_out_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_322 = _T_4112 ? dat_out_mask_38 : dl_out_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_323 = _T_4112 ? dat_out_mask_39 : dl_out_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_324 = _T_4112 ? dat_out_mask_40 : dl_out_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_325 = _T_4112 ? dat_out_mask_41 : dl_out_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_326 = _T_4112 ? dat_out_mask_42 : dl_out_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_327 = _T_4112 ? dat_out_mask_43 : dl_out_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_328 = _T_4112 ? dat_out_mask_44 : dl_out_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_329 = _T_4112 ? dat_out_mask_45 : dl_out_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_330 = _T_4112 ? dat_out_mask_46 : dl_out_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_331 = _T_4112 ? dat_out_mask_47 : dl_out_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_332 = _T_4112 ? dat_out_mask_48 : dl_out_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_333 = _T_4112 ? dat_out_mask_49 : dl_out_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_334 = _T_4112 ? dat_out_mask_50 : dl_out_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_335 = _T_4112 ? dat_out_mask_51 : dl_out_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_336 = _T_4112 ? dat_out_mask_52 : dl_out_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_337 = _T_4112 ? dat_out_mask_53 : dl_out_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_338 = _T_4112 ? dat_out_mask_54 : dl_out_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_339 = _T_4112 ? dat_out_mask_55 : dl_out_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_340 = _T_4112 ? dat_out_mask_56 : dl_out_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_341 = _T_4112 ? dat_out_mask_57 : dl_out_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_342 = _T_4112 ? dat_out_mask_58 : dl_out_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_343 = _T_4112 ? dat_out_mask_59 : dl_out_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_344 = _T_4112 ? dat_out_mask_60 : dl_out_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_345 = _T_4112 ? dat_out_mask_61 : dl_out_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_346 = _T_4112 ? dat_out_mask_62 : dl_out_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_347 = _T_4112 ? dat_out_mask_63 : dl_out_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1179:33:@2643.4]
  assign _GEN_348 = dat_out_pvld ? dat_out_flag : dl_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1182:19:@2709.4]
  assign _T_4115 = ~ dl_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:27:@2906.4]
  assign sc2mac_dat_pd_w = _T_4115 ? 9'h0 : dl_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1196:26:@2907.4]
  assign _T_4124 = dl_out_pvld | dl_out_pvld_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 1200:85:@2914.4]
  assign _GEN_413 = _T_4124 ? sc2mac_dat_pd_w : _T_4126; // @[Reg.scala 20:19:@2916.4]
  assign _GEN_414 = _T_4124 ? sc2mac_dat_pd_w : _T_4130; // @[Reg.scala 20:19:@2922.4]
  assign _GEN_415 = _T_4124 ? dl_out_mask_0 : _T_4398_0; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_416 = _T_4124 ? dl_out_mask_1 : _T_4398_1; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_417 = _T_4124 ? dl_out_mask_2 : _T_4398_2; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_418 = _T_4124 ? dl_out_mask_3 : _T_4398_3; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_419 = _T_4124 ? dl_out_mask_4 : _T_4398_4; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_420 = _T_4124 ? dl_out_mask_5 : _T_4398_5; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_421 = _T_4124 ? dl_out_mask_6 : _T_4398_6; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_422 = _T_4124 ? dl_out_mask_7 : _T_4398_7; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_423 = _T_4124 ? dl_out_mask_8 : _T_4398_8; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_424 = _T_4124 ? dl_out_mask_9 : _T_4398_9; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_425 = _T_4124 ? dl_out_mask_10 : _T_4398_10; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_426 = _T_4124 ? dl_out_mask_11 : _T_4398_11; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_427 = _T_4124 ? dl_out_mask_12 : _T_4398_12; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_428 = _T_4124 ? dl_out_mask_13 : _T_4398_13; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_429 = _T_4124 ? dl_out_mask_14 : _T_4398_14; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_430 = _T_4124 ? dl_out_mask_15 : _T_4398_15; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_431 = _T_4124 ? dl_out_mask_16 : _T_4398_16; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_432 = _T_4124 ? dl_out_mask_17 : _T_4398_17; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_433 = _T_4124 ? dl_out_mask_18 : _T_4398_18; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_434 = _T_4124 ? dl_out_mask_19 : _T_4398_19; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_435 = _T_4124 ? dl_out_mask_20 : _T_4398_20; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_436 = _T_4124 ? dl_out_mask_21 : _T_4398_21; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_437 = _T_4124 ? dl_out_mask_22 : _T_4398_22; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_438 = _T_4124 ? dl_out_mask_23 : _T_4398_23; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_439 = _T_4124 ? dl_out_mask_24 : _T_4398_24; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_440 = _T_4124 ? dl_out_mask_25 : _T_4398_25; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_441 = _T_4124 ? dl_out_mask_26 : _T_4398_26; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_442 = _T_4124 ? dl_out_mask_27 : _T_4398_27; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_443 = _T_4124 ? dl_out_mask_28 : _T_4398_28; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_444 = _T_4124 ? dl_out_mask_29 : _T_4398_29; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_445 = _T_4124 ? dl_out_mask_30 : _T_4398_30; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_446 = _T_4124 ? dl_out_mask_31 : _T_4398_31; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_447 = _T_4124 ? dl_out_mask_32 : _T_4398_32; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_448 = _T_4124 ? dl_out_mask_33 : _T_4398_33; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_449 = _T_4124 ? dl_out_mask_34 : _T_4398_34; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_450 = _T_4124 ? dl_out_mask_35 : _T_4398_35; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_451 = _T_4124 ? dl_out_mask_36 : _T_4398_36; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_452 = _T_4124 ? dl_out_mask_37 : _T_4398_37; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_453 = _T_4124 ? dl_out_mask_38 : _T_4398_38; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_454 = _T_4124 ? dl_out_mask_39 : _T_4398_39; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_455 = _T_4124 ? dl_out_mask_40 : _T_4398_40; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_456 = _T_4124 ? dl_out_mask_41 : _T_4398_41; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_457 = _T_4124 ? dl_out_mask_42 : _T_4398_42; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_458 = _T_4124 ? dl_out_mask_43 : _T_4398_43; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_459 = _T_4124 ? dl_out_mask_44 : _T_4398_44; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_460 = _T_4124 ? dl_out_mask_45 : _T_4398_45; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_461 = _T_4124 ? dl_out_mask_46 : _T_4398_46; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_462 = _T_4124 ? dl_out_mask_47 : _T_4398_47; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_463 = _T_4124 ? dl_out_mask_48 : _T_4398_48; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_464 = _T_4124 ? dl_out_mask_49 : _T_4398_49; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_465 = _T_4124 ? dl_out_mask_50 : _T_4398_50; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_466 = _T_4124 ? dl_out_mask_51 : _T_4398_51; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_467 = _T_4124 ? dl_out_mask_52 : _T_4398_52; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_468 = _T_4124 ? dl_out_mask_53 : _T_4398_53; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_469 = _T_4124 ? dl_out_mask_54 : _T_4398_54; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_470 = _T_4124 ? dl_out_mask_55 : _T_4398_55; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_471 = _T_4124 ? dl_out_mask_56 : _T_4398_56; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_472 = _T_4124 ? dl_out_mask_57 : _T_4398_57; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_473 = _T_4124 ? dl_out_mask_58 : _T_4398_58; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_474 = _T_4124 ? dl_out_mask_59 : _T_4398_59; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_475 = _T_4124 ? dl_out_mask_60 : _T_4398_60; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_476 = _T_4124 ? dl_out_mask_61 : _T_4398_61; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_477 = _T_4124 ? dl_out_mask_62 : _T_4398_62; // @[Reg.scala 20:19:@2993.4]
  assign _GEN_478 = _T_4124 ? dl_out_mask_63 : _T_4398_63; // @[Reg.scala 20:19:@2993.4]
  assign _T_4601 = {_T_4398_7,_T_4398_6,_T_4398_5,_T_4398_4,_T_4398_3,_T_4398_2,_T_4398_1,_T_4398_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3065.4]
  assign _T_4609 = {_T_4398_15,_T_4398_14,_T_4398_13,_T_4398_12,_T_4398_11,_T_4398_10,_T_4398_9,_T_4398_8,_T_4601}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3073.4]
  assign _T_4616 = {_T_4398_23,_T_4398_22,_T_4398_21,_T_4398_20,_T_4398_19,_T_4398_18,_T_4398_17,_T_4398_16}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3080.4]
  assign _T_4625 = {_T_4398_31,_T_4398_30,_T_4398_29,_T_4398_28,_T_4398_27,_T_4398_26,_T_4398_25,_T_4398_24,_T_4616,_T_4609}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3089.4]
  assign _T_4632 = {_T_4398_39,_T_4398_38,_T_4398_37,_T_4398_36,_T_4398_35,_T_4398_34,_T_4398_33,_T_4398_32}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3096.4]
  assign _T_4640 = {_T_4398_47,_T_4398_46,_T_4398_45,_T_4398_44,_T_4398_43,_T_4398_42,_T_4398_41,_T_4398_40,_T_4632}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3104.4]
  assign _T_4647 = {_T_4398_55,_T_4398_54,_T_4398_53,_T_4398_52,_T_4398_51,_T_4398_50,_T_4398_49,_T_4398_48}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3111.4]
  assign _T_4656 = {_T_4398_63,_T_4398_62,_T_4398_61,_T_4398_60,_T_4398_59,_T_4398_58,_T_4398_57,_T_4398_56,_T_4647,_T_4640}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:127:@3120.4]
  assign _GEN_479 = _T_4124 ? dl_out_mask_0 : _T_4925_0; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_480 = _T_4124 ? dl_out_mask_1 : _T_4925_1; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_481 = _T_4124 ? dl_out_mask_2 : _T_4925_2; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_482 = _T_4124 ? dl_out_mask_3 : _T_4925_3; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_483 = _T_4124 ? dl_out_mask_4 : _T_4925_4; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_484 = _T_4124 ? dl_out_mask_5 : _T_4925_5; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_485 = _T_4124 ? dl_out_mask_6 : _T_4925_6; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_486 = _T_4124 ? dl_out_mask_7 : _T_4925_7; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_487 = _T_4124 ? dl_out_mask_8 : _T_4925_8; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_488 = _T_4124 ? dl_out_mask_9 : _T_4925_9; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_489 = _T_4124 ? dl_out_mask_10 : _T_4925_10; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_490 = _T_4124 ? dl_out_mask_11 : _T_4925_11; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_491 = _T_4124 ? dl_out_mask_12 : _T_4925_12; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_492 = _T_4124 ? dl_out_mask_13 : _T_4925_13; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_493 = _T_4124 ? dl_out_mask_14 : _T_4925_14; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_494 = _T_4124 ? dl_out_mask_15 : _T_4925_15; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_495 = _T_4124 ? dl_out_mask_16 : _T_4925_16; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_496 = _T_4124 ? dl_out_mask_17 : _T_4925_17; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_497 = _T_4124 ? dl_out_mask_18 : _T_4925_18; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_498 = _T_4124 ? dl_out_mask_19 : _T_4925_19; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_499 = _T_4124 ? dl_out_mask_20 : _T_4925_20; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_500 = _T_4124 ? dl_out_mask_21 : _T_4925_21; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_501 = _T_4124 ? dl_out_mask_22 : _T_4925_22; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_502 = _T_4124 ? dl_out_mask_23 : _T_4925_23; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_503 = _T_4124 ? dl_out_mask_24 : _T_4925_24; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_504 = _T_4124 ? dl_out_mask_25 : _T_4925_25; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_505 = _T_4124 ? dl_out_mask_26 : _T_4925_26; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_506 = _T_4124 ? dl_out_mask_27 : _T_4925_27; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_507 = _T_4124 ? dl_out_mask_28 : _T_4925_28; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_508 = _T_4124 ? dl_out_mask_29 : _T_4925_29; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_509 = _T_4124 ? dl_out_mask_30 : _T_4925_30; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_510 = _T_4124 ? dl_out_mask_31 : _T_4925_31; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_511 = _T_4124 ? dl_out_mask_32 : _T_4925_32; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_512 = _T_4124 ? dl_out_mask_33 : _T_4925_33; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_513 = _T_4124 ? dl_out_mask_34 : _T_4925_34; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_514 = _T_4124 ? dl_out_mask_35 : _T_4925_35; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_515 = _T_4124 ? dl_out_mask_36 : _T_4925_36; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_516 = _T_4124 ? dl_out_mask_37 : _T_4925_37; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_517 = _T_4124 ? dl_out_mask_38 : _T_4925_38; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_518 = _T_4124 ? dl_out_mask_39 : _T_4925_39; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_519 = _T_4124 ? dl_out_mask_40 : _T_4925_40; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_520 = _T_4124 ? dl_out_mask_41 : _T_4925_41; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_521 = _T_4124 ? dl_out_mask_42 : _T_4925_42; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_522 = _T_4124 ? dl_out_mask_43 : _T_4925_43; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_523 = _T_4124 ? dl_out_mask_44 : _T_4925_44; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_524 = _T_4124 ? dl_out_mask_45 : _T_4925_45; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_525 = _T_4124 ? dl_out_mask_46 : _T_4925_46; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_526 = _T_4124 ? dl_out_mask_47 : _T_4925_47; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_527 = _T_4124 ? dl_out_mask_48 : _T_4925_48; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_528 = _T_4124 ? dl_out_mask_49 : _T_4925_49; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_529 = _T_4124 ? dl_out_mask_50 : _T_4925_50; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_530 = _T_4124 ? dl_out_mask_51 : _T_4925_51; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_531 = _T_4124 ? dl_out_mask_52 : _T_4925_52; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_532 = _T_4124 ? dl_out_mask_53 : _T_4925_53; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_533 = _T_4124 ? dl_out_mask_54 : _T_4925_54; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_534 = _T_4124 ? dl_out_mask_55 : _T_4925_55; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_535 = _T_4124 ? dl_out_mask_56 : _T_4925_56; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_536 = _T_4124 ? dl_out_mask_57 : _T_4925_57; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_537 = _T_4124 ? dl_out_mask_58 : _T_4925_58; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_538 = _T_4124 ? dl_out_mask_59 : _T_4925_59; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_539 = _T_4124 ? dl_out_mask_60 : _T_4925_60; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_540 = _T_4124 ? dl_out_mask_61 : _T_4925_61; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_541 = _T_4124 ? dl_out_mask_62 : _T_4925_62; // @[Reg.scala 20:19:@3190.4]
  assign _GEN_542 = _T_4124 ? dl_out_mask_63 : _T_4925_63; // @[Reg.scala 20:19:@3190.4]
  assign _T_5128 = {_T_4925_7,_T_4925_6,_T_4925_5,_T_4925_4,_T_4925_3,_T_4925_2,_T_4925_1,_T_4925_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3262.4]
  assign _T_5136 = {_T_4925_15,_T_4925_14,_T_4925_13,_T_4925_12,_T_4925_11,_T_4925_10,_T_4925_9,_T_4925_8,_T_5128}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3270.4]
  assign _T_5143 = {_T_4925_23,_T_4925_22,_T_4925_21,_T_4925_20,_T_4925_19,_T_4925_18,_T_4925_17,_T_4925_16}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3277.4]
  assign _T_5152 = {_T_4925_31,_T_4925_30,_T_4925_29,_T_4925_28,_T_4925_27,_T_4925_26,_T_4925_25,_T_4925_24,_T_5143,_T_5136}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3286.4]
  assign _T_5159 = {_T_4925_39,_T_4925_38,_T_4925_37,_T_4925_36,_T_4925_35,_T_4925_34,_T_4925_33,_T_4925_32}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3293.4]
  assign _T_5167 = {_T_4925_47,_T_4925_46,_T_4925_45,_T_4925_44,_T_4925_43,_T_4925_42,_T_4925_41,_T_4925_40,_T_5159}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3301.4]
  assign _T_5174 = {_T_4925_55,_T_4925_54,_T_4925_53,_T_4925_52,_T_4925_51,_T_4925_50,_T_4925_49,_T_4925_48}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3308.4]
  assign _T_5183 = {_T_4925_63,_T_4925_62,_T_4925_61,_T_4925_60,_T_4925_59,_T_4925_58,_T_4925_57,_T_4925_56,_T_5174,_T_5167}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:127:@3317.4]
  assign sc2cdma_dat_updt = _T_773; // @[NV_NVDLA_CSC_dl_for_check.scala 332:21:@325.4]
  assign sc2cdma_dat_entries = _T_779; // @[NV_NVDLA_CSC_dl_for_check.scala 334:24:@335.4]
  assign sc2cdma_dat_slices = _T_776; // @[NV_NVDLA_CSC_dl_for_check.scala 333:23:@330.4]
  assign sc2buf_dat_rd_en = sc2buf_dat_rd_en_out; // @[NV_NVDLA_CSC_dl_for_check.scala 749:29:@920.4]
  assign sc2buf_dat_rd_addr = sc2buf_dat_rd_addr_out[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 750:28:@921.4]
  assign sc2mac_dat_a_pvld = _T_4119; // @[NV_NVDLA_CSC_dl_for_check.scala 1198:23:@2910.4]
  assign sc2mac_dat_a_mask = {_T_4656,_T_4625}; // @[NV_NVDLA_CSC_dl_for_check.scala 1202:27:@3122.4]
  assign sc2mac_dat_a_data0 = _T_5186; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3324.4]
  assign sc2mac_dat_a_data1 = _T_5190; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3334.4]
  assign sc2mac_dat_a_data2 = _T_5194; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3344.4]
  assign sc2mac_dat_a_data3 = _T_5198; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3354.4]
  assign sc2mac_dat_a_data4 = _T_5202; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3364.4]
  assign sc2mac_dat_a_data5 = _T_5206; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3374.4]
  assign sc2mac_dat_a_data6 = _T_5210; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3384.4]
  assign sc2mac_dat_a_data7 = _T_5214; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3394.4]
  assign sc2mac_dat_a_data8 = _T_5218; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3404.4]
  assign sc2mac_dat_a_data9 = _T_5222; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3414.4]
  assign sc2mac_dat_a_data10 = _T_5226; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3424.4]
  assign sc2mac_dat_a_data11 = _T_5230; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3434.4]
  assign sc2mac_dat_a_data12 = _T_5234; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3444.4]
  assign sc2mac_dat_a_data13 = _T_5238; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3454.4]
  assign sc2mac_dat_a_data14 = _T_5242; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3464.4]
  assign sc2mac_dat_a_data15 = _T_5246; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3474.4]
  assign sc2mac_dat_a_data16 = _T_5250; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3484.4]
  assign sc2mac_dat_a_data17 = _T_5254; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3494.4]
  assign sc2mac_dat_a_data18 = _T_5258; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3504.4]
  assign sc2mac_dat_a_data19 = _T_5262; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3514.4]
  assign sc2mac_dat_a_data20 = _T_5266; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3524.4]
  assign sc2mac_dat_a_data21 = _T_5270; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3534.4]
  assign sc2mac_dat_a_data22 = _T_5274; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3544.4]
  assign sc2mac_dat_a_data23 = _T_5278; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3554.4]
  assign sc2mac_dat_a_data24 = _T_5282; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3564.4]
  assign sc2mac_dat_a_data25 = _T_5286; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3574.4]
  assign sc2mac_dat_a_data26 = _T_5290; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3584.4]
  assign sc2mac_dat_a_data27 = _T_5294; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3594.4]
  assign sc2mac_dat_a_data28 = _T_5298; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3604.4]
  assign sc2mac_dat_a_data29 = _T_5302; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3614.4]
  assign sc2mac_dat_a_data30 = _T_5306; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3624.4]
  assign sc2mac_dat_a_data31 = _T_5310; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3634.4]
  assign sc2mac_dat_a_data32 = _T_5314; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3644.4]
  assign sc2mac_dat_a_data33 = _T_5318; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3654.4]
  assign sc2mac_dat_a_data34 = _T_5322; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3664.4]
  assign sc2mac_dat_a_data35 = _T_5326; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3674.4]
  assign sc2mac_dat_a_data36 = _T_5330; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3684.4]
  assign sc2mac_dat_a_data37 = _T_5334; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3694.4]
  assign sc2mac_dat_a_data38 = _T_5338; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3704.4]
  assign sc2mac_dat_a_data39 = _T_5342; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3714.4]
  assign sc2mac_dat_a_data40 = _T_5346; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3724.4]
  assign sc2mac_dat_a_data41 = _T_5350; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3734.4]
  assign sc2mac_dat_a_data42 = _T_5354; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3744.4]
  assign sc2mac_dat_a_data43 = _T_5358; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3754.4]
  assign sc2mac_dat_a_data44 = _T_5362; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3764.4]
  assign sc2mac_dat_a_data45 = _T_5366; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3774.4]
  assign sc2mac_dat_a_data46 = _T_5370; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3784.4]
  assign sc2mac_dat_a_data47 = _T_5374; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3794.4]
  assign sc2mac_dat_a_data48 = _T_5378; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3804.4]
  assign sc2mac_dat_a_data49 = _T_5382; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3814.4]
  assign sc2mac_dat_a_data50 = _T_5386; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3824.4]
  assign sc2mac_dat_a_data51 = _T_5390; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3834.4]
  assign sc2mac_dat_a_data52 = _T_5394; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3844.4]
  assign sc2mac_dat_a_data53 = _T_5398; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3854.4]
  assign sc2mac_dat_a_data54 = _T_5402; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3864.4]
  assign sc2mac_dat_a_data55 = _T_5406; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3874.4]
  assign sc2mac_dat_a_data56 = _T_5410; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3884.4]
  assign sc2mac_dat_a_data57 = _T_5414; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3894.4]
  assign sc2mac_dat_a_data58 = _T_5418; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3904.4]
  assign sc2mac_dat_a_data59 = _T_5422; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3914.4]
  assign sc2mac_dat_a_data60 = _T_5426; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3924.4]
  assign sc2mac_dat_a_data61 = _T_5430; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3934.4]
  assign sc2mac_dat_a_data62 = _T_5434; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3944.4]
  assign sc2mac_dat_a_data63 = _T_5438; // @[NV_NVDLA_CSC_dl_for_check.scala 1205:34:@3954.4]
  assign sc2mac_dat_a_pd = _T_4126; // @[NV_NVDLA_CSC_dl_for_check.scala 1200:25:@2919.4]
  assign sc2mac_dat_b_pvld = _T_4122; // @[NV_NVDLA_CSC_dl_for_check.scala 1199:23:@2913.4]
  assign sc2mac_dat_b_mask = {_T_5183,_T_5152}; // @[NV_NVDLA_CSC_dl_for_check.scala 1203:27:@3319.4]
  assign sc2mac_dat_b_data0 = _T_5188; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3329.4]
  assign sc2mac_dat_b_data1 = _T_5192; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3339.4]
  assign sc2mac_dat_b_data2 = _T_5196; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3349.4]
  assign sc2mac_dat_b_data3 = _T_5200; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3359.4]
  assign sc2mac_dat_b_data4 = _T_5204; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3369.4]
  assign sc2mac_dat_b_data5 = _T_5208; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3379.4]
  assign sc2mac_dat_b_data6 = _T_5212; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3389.4]
  assign sc2mac_dat_b_data7 = _T_5216; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3399.4]
  assign sc2mac_dat_b_data8 = _T_5220; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3409.4]
  assign sc2mac_dat_b_data9 = _T_5224; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3419.4]
  assign sc2mac_dat_b_data10 = _T_5228; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3429.4]
  assign sc2mac_dat_b_data11 = _T_5232; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3439.4]
  assign sc2mac_dat_b_data12 = _T_5236; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3449.4]
  assign sc2mac_dat_b_data13 = _T_5240; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3459.4]
  assign sc2mac_dat_b_data14 = _T_5244; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3469.4]
  assign sc2mac_dat_b_data15 = _T_5248; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3479.4]
  assign sc2mac_dat_b_data16 = _T_5252; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3489.4]
  assign sc2mac_dat_b_data17 = _T_5256; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3499.4]
  assign sc2mac_dat_b_data18 = _T_5260; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3509.4]
  assign sc2mac_dat_b_data19 = _T_5264; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3519.4]
  assign sc2mac_dat_b_data20 = _T_5268; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3529.4]
  assign sc2mac_dat_b_data21 = _T_5272; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3539.4]
  assign sc2mac_dat_b_data22 = _T_5276; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3549.4]
  assign sc2mac_dat_b_data23 = _T_5280; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3559.4]
  assign sc2mac_dat_b_data24 = _T_5284; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3569.4]
  assign sc2mac_dat_b_data25 = _T_5288; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3579.4]
  assign sc2mac_dat_b_data26 = _T_5292; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3589.4]
  assign sc2mac_dat_b_data27 = _T_5296; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3599.4]
  assign sc2mac_dat_b_data28 = _T_5300; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3609.4]
  assign sc2mac_dat_b_data29 = _T_5304; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3619.4]
  assign sc2mac_dat_b_data30 = _T_5308; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3629.4]
  assign sc2mac_dat_b_data31 = _T_5312; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3639.4]
  assign sc2mac_dat_b_data32 = _T_5316; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3649.4]
  assign sc2mac_dat_b_data33 = _T_5320; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3659.4]
  assign sc2mac_dat_b_data34 = _T_5324; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3669.4]
  assign sc2mac_dat_b_data35 = _T_5328; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3679.4]
  assign sc2mac_dat_b_data36 = _T_5332; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3689.4]
  assign sc2mac_dat_b_data37 = _T_5336; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3699.4]
  assign sc2mac_dat_b_data38 = _T_5340; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3709.4]
  assign sc2mac_dat_b_data39 = _T_5344; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3719.4]
  assign sc2mac_dat_b_data40 = _T_5348; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3729.4]
  assign sc2mac_dat_b_data41 = _T_5352; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3739.4]
  assign sc2mac_dat_b_data42 = _T_5356; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3749.4]
  assign sc2mac_dat_b_data43 = _T_5360; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3759.4]
  assign sc2mac_dat_b_data44 = _T_5364; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3769.4]
  assign sc2mac_dat_b_data45 = _T_5368; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3779.4]
  assign sc2mac_dat_b_data46 = _T_5372; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3789.4]
  assign sc2mac_dat_b_data47 = _T_5376; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3799.4]
  assign sc2mac_dat_b_data48 = _T_5380; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3809.4]
  assign sc2mac_dat_b_data49 = _T_5384; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3819.4]
  assign sc2mac_dat_b_data50 = _T_5388; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3829.4]
  assign sc2mac_dat_b_data51 = _T_5392; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3839.4]
  assign sc2mac_dat_b_data52 = _T_5396; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3849.4]
  assign sc2mac_dat_b_data53 = _T_5400; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3859.4]
  assign sc2mac_dat_b_data54 = _T_5404; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3869.4]
  assign sc2mac_dat_b_data55 = _T_5408; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3879.4]
  assign sc2mac_dat_b_data56 = _T_5412; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3889.4]
  assign sc2mac_dat_b_data57 = _T_5416; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3899.4]
  assign sc2mac_dat_b_data58 = _T_5420; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3909.4]
  assign sc2mac_dat_b_data59 = _T_5424; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3919.4]
  assign sc2mac_dat_b_data60 = _T_5428; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3929.4]
  assign sc2mac_dat_b_data61 = _T_5432; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3939.4]
  assign sc2mac_dat_b_data62 = _T_5436; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3949.4]
  assign sc2mac_dat_b_data63 = _T_5440; // @[NV_NVDLA_CSC_dl_for_check.scala 1206:34:@3959.4]
  assign sc2mac_dat_b_pd = _T_4130; // @[NV_NVDLA_CSC_dl_for_check.scala 1201:25:@2925.4]
  assign slcg_wg_en = 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 273:15:@242.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  layer_st_d1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_batch = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rls_slices = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  h_offset_slice = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  entries = _RAND_4[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  entries_batch = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  dataout_width_cmp = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rls_entries = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  h_bias_0_stride = _RAND_8[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  h_bias_1_stride = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  slice_left = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {2{`RANDOM}};
  is_img_d1 = _RAND_11[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  data_bank = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  datain_width = _RAND_13[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  datain_width_cmp = _RAND_14[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  datain_height_cmp = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  datain_channel_cmp = _RAND_16[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  sub_h_total_g0 = _RAND_17[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sub_h_total_g1 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  sub_h_total_g3 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  sub_h_total_g4 = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  sub_h_total_g5 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  sub_h_total_g6 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sub_h_total_g8 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sub_h_total_g9 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sub_h_total_g11 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sub_h_cmp_g0 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sub_h_cmp_g1 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  conv_x_stride = _RAND_28[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  conv_y_stride = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  batch_cmp = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  pixel_x_init = _RAND_31[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  pixel_x_init_offset = _RAND_32[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  pixel_x_add = _RAND_33[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  pixel_x_byte_stride = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  pixel_ch_stride = _RAND_35[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  x_dilate = _RAND_36[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  y_dilate = _RAND_37[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  pad_value = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  entries_cmp = _RAND_39[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  h_bias_2_stride = _RAND_40[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  h_bias_3_stride = _RAND_41[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  last_slices = _RAND_42[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  last_entries = _RAND_43[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  dat_entry_st = _RAND_44[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  dat_rsp_l3_pvld = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  dat_rsp_l1_pvld = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  dat_rsp_l0_pvld = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_1617 = _RAND_48[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_1611 = _RAND_49[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1608 = _RAND_50[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_773 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_776 = _RAND_52[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_779 = _RAND_53[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_784 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_787 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_790 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_793 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  dl_in_pvld = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_817 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_820 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_823 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_826 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_831 = _RAND_63[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_834 = _RAND_64[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_837 = _RAND_65[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_840 = _RAND_66[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  batch_cnt = _RAND_67[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  sub_h_cnt = _RAND_68[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  stripe_cnt = _RAND_69[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  dat_exec_valid_d1 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  dat_pipe_local_valid = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  dat_pipe_valid_d1 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  dat_req_bytes_d1 = _RAND_73[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  dataout_w_cnt = _RAND_74[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  dataout_w_ori = _RAND_75[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  datain_c_cnt = _RAND_76[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  datain_w_cnt = _RAND_77[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  datain_w_ori = _RAND_78[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  pixel_w_cnt = _RAND_79[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  pixel_w_ori = _RAND_80[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  pixel_w_ch_ori = _RAND_81[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  channel_op_cnt = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  pixel_force_clr_d1 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  pixel_force_fetch_d1 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  datain_h_cnt = _RAND_85[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  datain_h_ori = _RAND_86[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  dat_req_valid_d1 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  dat_req_sub_w_d1 = _RAND_88[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  dat_req_sub_h_d1 = _RAND_89[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  dat_req_sub_c_d1 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  dat_req_ch_end_d1 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  dat_req_dummy_d1 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  dat_req_cur_sub_h_d1 = _RAND_93[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dat_req_sub_w_st_d1 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dat_req_flag_d1 = _RAND_95[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dat_req_rls_d1 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  c_bias = _RAND_97[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  c_bias_d1 = _RAND_98[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  h_bias_0_d1 = _RAND_99[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  h_bias_1_d1 = _RAND_100[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  h_bias_2_d1 = _RAND_101[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  h_bias_3_d1 = _RAND_102[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  w_bias_d1 = _RAND_103[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  dat_req_sub_h_addr_0 = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  dat_req_sub_h_addr_1 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  dat_req_sub_h_addr_2 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  sc2buf_dat_rd_en_out = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  sc2buf_dat_rd_addr_out = _RAND_108[17:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  dat_req_pipe_pvld = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  dat_req_pipe_sub_w = _RAND_110[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  dat_req_pipe_sub_h = _RAND_111[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  dat_req_pipe_sub_c = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  dat_req_pipe_ch_end = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  dat_req_pipe_bytes = _RAND_114[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  dat_req_pipe_dummy = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  dat_req_pipe_cur_sub_h = _RAND_116[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  dat_req_pipe_sub_w_st = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  dat_req_pipe_rls = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  dat_req_pipe_flag = _RAND_119[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_1389 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_1392 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_1395 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_1398 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_1401 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  dat_rsp_pipe_pvld = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_1408 = _RAND_126[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_1411 = _RAND_127[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_1414 = _RAND_128[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_1417 = _RAND_129[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1420 = _RAND_130[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  dat_rsp_pipe_pd = _RAND_131[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  dat_l0c0_dummy = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  dat_l0c1_dummy = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {16{`RANDOM}};
  dat_l0c0 = _RAND_134[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {16{`RANDOM}};
  dat_l0c1 = _RAND_135[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  rsp_sft_cnt_l0 = _RAND_136[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  rsp_sft_cnt_l1 = _RAND_137[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  rsp_sft_cnt_l2 = _RAND_138[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  rsp_sft_cnt_l3 = _RAND_139[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  rsp_sft_cnt_l0_ori = _RAND_140[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  rsp_sft_cnt_l1_ori = _RAND_141[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  rsp_sft_cnt_l2_ori = _RAND_142[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  rsp_sft_cnt_l3_ori = _RAND_143[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  dat_rsp_l2_pvld = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_1614 = _RAND_145[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {8{`RANDOM}};
  dat_rsp_l0_sft_d1 = _RAND_146[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {4{`RANDOM}};
  dat_rsp_l0_sft_d2 = _RAND_147[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {4{`RANDOM}};
  dat_rsp_l0_sft_d3 = _RAND_148[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {4{`RANDOM}};
  dat_rsp_l1_sft_d2 = _RAND_149[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {4{`RANDOM}};
  dat_rsp_l1_sft_d3 = _RAND_150[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {4{`RANDOM}};
  dat_rsp_l2_sft_d3 = _RAND_151[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  dat_out_pvld = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  dat_out_flag = _RAND_153[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  dat_out_bypass_mask_0 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  dat_out_bypass_mask_1 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  dat_out_bypass_mask_2 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  dat_out_bypass_mask_3 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  dat_out_bypass_mask_4 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  dat_out_bypass_mask_5 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  dat_out_bypass_mask_6 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  dat_out_bypass_mask_7 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  dat_out_bypass_mask_8 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  dat_out_bypass_mask_9 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  dat_out_bypass_mask_10 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  dat_out_bypass_mask_11 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  dat_out_bypass_mask_12 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  dat_out_bypass_mask_13 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  dat_out_bypass_mask_14 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  dat_out_bypass_mask_15 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  dat_out_bypass_mask_16 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  dat_out_bypass_mask_17 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  dat_out_bypass_mask_18 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  dat_out_bypass_mask_19 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  dat_out_bypass_mask_20 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  dat_out_bypass_mask_21 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  dat_out_bypass_mask_22 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  dat_out_bypass_mask_23 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  dat_out_bypass_mask_24 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  dat_out_bypass_mask_25 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  dat_out_bypass_mask_26 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  dat_out_bypass_mask_27 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  dat_out_bypass_mask_28 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  dat_out_bypass_mask_29 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  dat_out_bypass_mask_30 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  dat_out_bypass_mask_31 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  dat_out_bypass_mask_32 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  dat_out_bypass_mask_33 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  dat_out_bypass_mask_34 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  dat_out_bypass_mask_35 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  dat_out_bypass_mask_36 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  dat_out_bypass_mask_37 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  dat_out_bypass_mask_38 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  dat_out_bypass_mask_39 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  dat_out_bypass_mask_40 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  dat_out_bypass_mask_41 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  dat_out_bypass_mask_42 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  dat_out_bypass_mask_43 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  dat_out_bypass_mask_44 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  dat_out_bypass_mask_45 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  dat_out_bypass_mask_46 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  dat_out_bypass_mask_47 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  dat_out_bypass_mask_48 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  dat_out_bypass_mask_49 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  dat_out_bypass_mask_50 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  dat_out_bypass_mask_51 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  dat_out_bypass_mask_52 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  dat_out_bypass_mask_53 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  dat_out_bypass_mask_54 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  dat_out_bypass_mask_55 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  dat_out_bypass_mask_56 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  dat_out_bypass_mask_57 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  dat_out_bypass_mask_58 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  dat_out_bypass_mask_59 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  dat_out_bypass_mask_60 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  dat_out_bypass_mask_61 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  dat_out_bypass_mask_62 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  dat_out_bypass_mask_63 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  dat_out_bypass_data_0 = _RAND_218[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  dat_out_bypass_data_1 = _RAND_219[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  dat_out_bypass_data_2 = _RAND_220[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  dat_out_bypass_data_3 = _RAND_221[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  dat_out_bypass_data_4 = _RAND_222[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  dat_out_bypass_data_5 = _RAND_223[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  dat_out_bypass_data_6 = _RAND_224[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  dat_out_bypass_data_7 = _RAND_225[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  dat_out_bypass_data_8 = _RAND_226[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  dat_out_bypass_data_9 = _RAND_227[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  dat_out_bypass_data_10 = _RAND_228[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  dat_out_bypass_data_11 = _RAND_229[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  dat_out_bypass_data_12 = _RAND_230[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  dat_out_bypass_data_13 = _RAND_231[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  dat_out_bypass_data_14 = _RAND_232[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  dat_out_bypass_data_15 = _RAND_233[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  dat_out_bypass_data_16 = _RAND_234[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  dat_out_bypass_data_17 = _RAND_235[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  dat_out_bypass_data_18 = _RAND_236[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  dat_out_bypass_data_19 = _RAND_237[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  dat_out_bypass_data_20 = _RAND_238[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  dat_out_bypass_data_21 = _RAND_239[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  dat_out_bypass_data_22 = _RAND_240[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  dat_out_bypass_data_23 = _RAND_241[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  dat_out_bypass_data_24 = _RAND_242[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  dat_out_bypass_data_25 = _RAND_243[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  dat_out_bypass_data_26 = _RAND_244[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  dat_out_bypass_data_27 = _RAND_245[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  dat_out_bypass_data_28 = _RAND_246[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  dat_out_bypass_data_29 = _RAND_247[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  dat_out_bypass_data_30 = _RAND_248[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  dat_out_bypass_data_31 = _RAND_249[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  dat_out_bypass_data_32 = _RAND_250[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  dat_out_bypass_data_33 = _RAND_251[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  dat_out_bypass_data_34 = _RAND_252[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  dat_out_bypass_data_35 = _RAND_253[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  dat_out_bypass_data_36 = _RAND_254[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  dat_out_bypass_data_37 = _RAND_255[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  dat_out_bypass_data_38 = _RAND_256[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  dat_out_bypass_data_39 = _RAND_257[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  dat_out_bypass_data_40 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  dat_out_bypass_data_41 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  dat_out_bypass_data_42 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  dat_out_bypass_data_43 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  dat_out_bypass_data_44 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  dat_out_bypass_data_45 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  dat_out_bypass_data_46 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  dat_out_bypass_data_47 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  dat_out_bypass_data_48 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  dat_out_bypass_data_49 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  dat_out_bypass_data_50 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  dat_out_bypass_data_51 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  dat_out_bypass_data_52 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  dat_out_bypass_data_53 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  dat_out_bypass_data_54 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  dat_out_bypass_data_55 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  dat_out_bypass_data_56 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  dat_out_bypass_data_57 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  dat_out_bypass_data_58 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  dat_out_bypass_data_59 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  dat_out_bypass_data_60 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  dat_out_bypass_data_61 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  dat_out_bypass_data_62 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  dat_out_bypass_data_63 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  dl_out_pvld = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  dl_out_mask_0 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  dl_out_mask_1 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  dl_out_mask_2 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  dl_out_mask_3 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  dl_out_mask_4 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  dl_out_mask_5 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  dl_out_mask_6 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  dl_out_mask_7 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  dl_out_mask_8 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  dl_out_mask_9 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  dl_out_mask_10 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  dl_out_mask_11 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  dl_out_mask_12 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  dl_out_mask_13 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  dl_out_mask_14 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  dl_out_mask_15 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  dl_out_mask_16 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  dl_out_mask_17 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  dl_out_mask_18 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  dl_out_mask_19 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  dl_out_mask_20 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  dl_out_mask_21 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  dl_out_mask_22 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  dl_out_mask_23 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  dl_out_mask_24 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  dl_out_mask_25 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  dl_out_mask_26 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  dl_out_mask_27 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  dl_out_mask_28 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  dl_out_mask_29 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  dl_out_mask_30 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  dl_out_mask_31 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  dl_out_mask_32 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  dl_out_mask_33 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  dl_out_mask_34 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  dl_out_mask_35 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  dl_out_mask_36 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  dl_out_mask_37 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  dl_out_mask_38 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  dl_out_mask_39 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  dl_out_mask_40 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  dl_out_mask_41 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  dl_out_mask_42 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  dl_out_mask_43 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  dl_out_mask_44 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  dl_out_mask_45 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  dl_out_mask_46 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  dl_out_mask_47 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  dl_out_mask_48 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  dl_out_mask_49 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  dl_out_mask_50 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  dl_out_mask_51 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  dl_out_mask_52 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  dl_out_mask_53 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  dl_out_mask_54 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  dl_out_mask_55 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  dl_out_mask_56 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  dl_out_mask_57 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  dl_out_mask_58 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  dl_out_mask_59 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  dl_out_mask_60 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  dl_out_mask_61 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  dl_out_mask_62 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  dl_out_mask_63 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  dl_out_flag = _RAND_347[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  dl_out_data_0 = _RAND_348[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  dl_out_data_1 = _RAND_349[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  dl_out_data_2 = _RAND_350[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  dl_out_data_3 = _RAND_351[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  dl_out_data_4 = _RAND_352[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  dl_out_data_5 = _RAND_353[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  dl_out_data_6 = _RAND_354[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  dl_out_data_7 = _RAND_355[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  dl_out_data_8 = _RAND_356[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  dl_out_data_9 = _RAND_357[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  dl_out_data_10 = _RAND_358[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  dl_out_data_11 = _RAND_359[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  dl_out_data_12 = _RAND_360[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  dl_out_data_13 = _RAND_361[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  dl_out_data_14 = _RAND_362[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  dl_out_data_15 = _RAND_363[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  dl_out_data_16 = _RAND_364[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  dl_out_data_17 = _RAND_365[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  dl_out_data_18 = _RAND_366[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  dl_out_data_19 = _RAND_367[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  dl_out_data_20 = _RAND_368[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  dl_out_data_21 = _RAND_369[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  dl_out_data_22 = _RAND_370[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  dl_out_data_23 = _RAND_371[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  dl_out_data_24 = _RAND_372[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  dl_out_data_25 = _RAND_373[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  dl_out_data_26 = _RAND_374[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  dl_out_data_27 = _RAND_375[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  dl_out_data_28 = _RAND_376[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  dl_out_data_29 = _RAND_377[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  dl_out_data_30 = _RAND_378[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  dl_out_data_31 = _RAND_379[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  dl_out_data_32 = _RAND_380[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  dl_out_data_33 = _RAND_381[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  dl_out_data_34 = _RAND_382[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  dl_out_data_35 = _RAND_383[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  dl_out_data_36 = _RAND_384[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  dl_out_data_37 = _RAND_385[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  dl_out_data_38 = _RAND_386[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  dl_out_data_39 = _RAND_387[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  dl_out_data_40 = _RAND_388[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  dl_out_data_41 = _RAND_389[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  dl_out_data_42 = _RAND_390[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  dl_out_data_43 = _RAND_391[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  dl_out_data_44 = _RAND_392[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  dl_out_data_45 = _RAND_393[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  dl_out_data_46 = _RAND_394[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  dl_out_data_47 = _RAND_395[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  dl_out_data_48 = _RAND_396[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  dl_out_data_49 = _RAND_397[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  dl_out_data_50 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  dl_out_data_51 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  dl_out_data_52 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  dl_out_data_53 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  dl_out_data_54 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  dl_out_data_55 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  dl_out_data_56 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  dl_out_data_57 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  dl_out_data_58 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  dl_out_data_59 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  dl_out_data_60 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  dl_out_data_61 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  dl_out_data_62 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  dl_out_data_63 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  dl_out_pvld_d1 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_4119 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_4122 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_4126 = _RAND_415[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_4130 = _RAND_416[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_4398_0 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_4398_1 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_4398_2 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_4398_3 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_4398_4 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_4398_5 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_4398_6 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_4398_7 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_4398_8 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_4398_9 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_4398_10 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_4398_11 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_4398_12 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_4398_13 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_4398_14 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_4398_15 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_4398_16 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_4398_17 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_4398_18 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_4398_19 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_4398_20 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_4398_21 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_4398_22 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_4398_23 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_4398_24 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_4398_25 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_4398_26 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_4398_27 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_4398_28 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_4398_29 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_4398_30 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_4398_31 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_4398_32 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_4398_33 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_4398_34 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_4398_35 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_4398_36 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_4398_37 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_4398_38 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_4398_39 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_4398_40 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_4398_41 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_4398_42 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_4398_43 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_4398_44 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_4398_45 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_4398_46 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_4398_47 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_4398_48 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_4398_49 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_4398_50 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_4398_51 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_4398_52 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_4398_53 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_4398_54 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_4398_55 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_4398_56 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_4398_57 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_4398_58 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_4398_59 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_4398_60 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_4398_61 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_4398_62 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_4398_63 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_4925_0 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_4925_1 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_4925_2 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_4925_3 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_4925_4 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_4925_5 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_4925_6 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_4925_7 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_4925_8 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_4925_9 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_4925_10 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_4925_11 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_4925_12 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_4925_13 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_4925_14 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_4925_15 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_4925_16 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_4925_17 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_4925_18 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_4925_19 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_4925_20 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_4925_21 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_4925_22 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_4925_23 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_4925_24 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_4925_25 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_4925_26 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_4925_27 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_4925_28 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_4925_29 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_4925_30 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_4925_31 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_4925_32 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_4925_33 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_4925_34 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_4925_35 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_4925_36 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_4925_37 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_4925_38 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_4925_39 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_4925_40 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_4925_41 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_4925_42 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_4925_43 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_4925_44 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_4925_45 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_4925_46 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_4925_47 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_4925_48 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_4925_49 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_4925_50 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_4925_51 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_4925_52 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_4925_53 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_4925_54 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_4925_55 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_4925_56 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_4925_57 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_4925_58 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_4925_59 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_4925_60 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_4925_61 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_4925_62 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_4925_63 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5186 = _RAND_545[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5188 = _RAND_546[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5190 = _RAND_547[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5192 = _RAND_548[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5194 = _RAND_549[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_5196 = _RAND_550[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_5198 = _RAND_551[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_5200 = _RAND_552[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_5202 = _RAND_553[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_5204 = _RAND_554[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_5206 = _RAND_555[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_5208 = _RAND_556[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_5210 = _RAND_557[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_5212 = _RAND_558[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_5214 = _RAND_559[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_5216 = _RAND_560[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_5218 = _RAND_561[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_5220 = _RAND_562[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_5222 = _RAND_563[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_5224 = _RAND_564[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_5226 = _RAND_565[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_5228 = _RAND_566[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_5230 = _RAND_567[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_5232 = _RAND_568[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_5234 = _RAND_569[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_5236 = _RAND_570[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_5238 = _RAND_571[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_5240 = _RAND_572[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_5242 = _RAND_573[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_5244 = _RAND_574[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_5246 = _RAND_575[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_5248 = _RAND_576[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_5250 = _RAND_577[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_5252 = _RAND_578[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_5254 = _RAND_579[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_5256 = _RAND_580[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_5258 = _RAND_581[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_5260 = _RAND_582[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_5262 = _RAND_583[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_5264 = _RAND_584[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_5266 = _RAND_585[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_5268 = _RAND_586[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_5270 = _RAND_587[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_5272 = _RAND_588[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_5274 = _RAND_589[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_5276 = _RAND_590[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_5278 = _RAND_591[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_5280 = _RAND_592[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_5282 = _RAND_593[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_5284 = _RAND_594[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_5286 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_5288 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_5290 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_5292 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_5294 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_5296 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_5298 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_5300 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_5302 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_5304 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_5306 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_5308 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_5310 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_5312 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_5314 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_5316 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_5318 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_5320 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_5322 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_5324 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_5326 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_5328 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_5330 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_5332 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_5334 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_5336 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_5338 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_5340 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_5342 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_5344 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_5346 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_5348 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_5350 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_5352 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_5354 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_5356 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_5358 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_5360 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_5362 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_5364 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_5366 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_5368 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_5370 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_5372 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_5374 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_5376 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_5378 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_5380 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_5382 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_5384 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_5386 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_5388 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_5390 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_5392 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_5394 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_5396 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_5398 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_5400 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_5402 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_5404 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_5406 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_5408 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_5410 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_5412 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_5414 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_5416 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_5418 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_5420 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_5422 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_5424 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_5426 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_5428 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_5430 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_5432 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_5434 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_5436 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_5438 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_5440 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge nvdla_core_clk) begin
    if (_T_337) begin
      layer_st_d1 <= 1'h0;
    end else begin
      layer_st_d1 <= layer_st;
    end
    if (_T_337) begin
      data_batch <= 6'h0;
    end else begin
      if (layer_st) begin
        data_batch <= 6'h1;
      end
    end
    if (_T_337) begin
      rls_slices <= 14'h0;
    end else begin
      if (layer_st) begin
        rls_slices <= {{1'd0}, rls_slices_w};
      end
    end
    if (_T_337) begin
      h_offset_slice <= 14'h0;
    end else begin
      if (layer_st) begin
        h_offset_slice <= {{2'd0}, h_offset_slice_w};
      end
    end
    if (_T_337) begin
      entries <= 15'h0;
    end else begin
      if (layer_st) begin
        entries <= entries_single_w;
      end
    end
    if (_T_337) begin
      entries_batch <= 15'h0;
    end else begin
      if (layer_st) begin
        entries_batch <= entries_batch_w;
      end
    end
    if (_T_337) begin
      dataout_width_cmp <= 13'h0;
    end else begin
      if (layer_st) begin
        dataout_width_cmp <= reg2dp_dataout_width;
      end
    end
    if (_T_337) begin
      rls_entries <= 15'h0;
    end else begin
      if (layer_st_d1) begin
        rls_entries <= slice_entries_w;
      end
    end
    if (_T_337) begin
      h_bias_0_stride <= 12'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_0_stride <= h_bias_0_stride_w;
      end
    end
    if (_T_337) begin
      h_bias_1_stride <= 12'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_1_stride <= h_bias_1_stride_w;
      end
    end
    if (_T_337) begin
      slice_left <= 14'h0;
    end else begin
      if (layer_st) begin
        if (reg2dp_skip_data_rls) begin
          slice_left <= _T_482;
        end else begin
          slice_left <= _T_484;
        end
      end
    end
    if (_T_337) begin
      is_img_d1 <= 34'h0;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          is_img_d1 <= 34'h3ffffffff;
        end else begin
          is_img_d1 <= 34'h0;
        end
      end
    end
    if (_T_337) begin
      data_bank <= 5'h0;
    end else begin
      if (layer_st) begin
        data_bank <= _T_673;
      end
    end
    if (_T_337) begin
      datain_width <= 14'h0;
    end else begin
      if (layer_st) begin
        datain_width <= _T_675;
      end
    end
    if (_T_337) begin
      datain_width_cmp <= 13'h0;
    end else begin
      if (layer_st) begin
        datain_width_cmp <= reg2dp_datain_width_ext;
      end
    end
    if (_T_337) begin
      datain_height_cmp <= 13'h0;
    end else begin
      if (layer_st) begin
        datain_height_cmp <= reg2dp_datain_height_ext;
      end
    end
    if (_T_337) begin
      datain_channel_cmp <= 11'h0;
    end else begin
      if (layer_st) begin
        datain_channel_cmp <= _T_682;
      end
    end
    if (_T_337) begin
      sub_h_total_g0 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g0 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g1 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g1 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g3 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g3 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g4 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g4 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g5 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g5 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g6 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g6 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g8 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g8 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g9 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g9 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_total_g11 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g11 <= sub_h_total_w;
      end
    end
    if (_T_337) begin
      sub_h_cmp_g0 <= 3'h1;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          sub_h_cmp_g0 <= sub_h_total_w;
        end else begin
          sub_h_cmp_g0 <= 3'h1;
        end
      end
    end
    if (_T_337) begin
      sub_h_cmp_g1 <= 3'h1;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          sub_h_cmp_g1 <= sub_h_total_w;
        end else begin
          sub_h_cmp_g1 <= 3'h1;
        end
      end
    end
    if (_T_337) begin
      conv_x_stride <= 4'h0;
    end else begin
      if (layer_st) begin
        conv_x_stride <= conv_x_stride_w;
      end
    end
    if (_T_337) begin
      conv_y_stride <= 4'h0;
    end else begin
      if (layer_st) begin
        conv_y_stride <= conv_y_stride_w;
      end
    end
    if (_T_337) begin
      batch_cmp <= 5'h0;
    end else begin
      if (layer_st) begin
        batch_cmp <= 5'h0;
      end
    end
    if (_T_337) begin
      pixel_x_init <= 7'h0;
    end else begin
      if (layer_st) begin
        if (_T_387) begin
          pixel_x_init <= _T_380;
        end else begin
          pixel_x_init <= {{1'd0}, _T_386};
        end
      end
    end
    if (_T_337) begin
      pixel_x_init_offset <= 7'h0;
    end else begin
      if (layer_st) begin
        pixel_x_init_offset <= pixel_x_init_offset_w;
      end
    end
    if (_T_337) begin
      pixel_x_add <= 8'h0;
    end else begin
      if (layer_st) begin
        if (_T_387) begin
          pixel_x_add <= _T_392;
        end else begin
          pixel_x_add <= {{1'd0}, _T_397};
        end
      end
    end
    if (_T_337) begin
      pixel_x_byte_stride <= 7'h0;
    end else begin
      if (layer_st) begin
        pixel_x_byte_stride <= {{1'd0}, pixel_x_stride_w};
      end
    end
    if (_T_337) begin
      pixel_ch_stride <= 12'h0;
    end else begin
      if (layer_st) begin
        pixel_ch_stride <= pixel_ch_stride_w;
      end
    end
    if (_T_337) begin
      x_dilate <= 6'h0;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          x_dilate <= 6'h1;
        end else begin
          x_dilate <= _T_403;
        end
      end
    end
    if (_T_337) begin
      y_dilate <= 6'h0;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          y_dilate <= 6'h1;
        end else begin
          y_dilate <= _T_406;
        end
      end
    end
    if (_T_337) begin
      pad_value <= 16'h0;
    end else begin
      if (layer_st) begin
        pad_value <= reg2dp_pad_value;
      end
    end
    if (_T_337) begin
      entries_cmp <= 15'h0;
    end else begin
      if (layer_st) begin
        entries_cmp <= _T_686;
      end
    end
    if (_T_337) begin
      h_bias_2_stride <= 15'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_2_stride <= entries;
      end
    end
    if (_T_337) begin
      h_bias_3_stride <= 15'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_3_stride <= entries;
      end
    end
    if (_T_337) begin
      last_slices <= 14'h0;
    end else begin
      if (is_sg_done) begin
        last_slices <= slice_left;
      end
    end
    if (_T_337) begin
      last_entries <= 15'h0;
    end else begin
      if (is_sg_done) begin
        last_entries <= slice_entries_w;
      end
    end
    if (_T_337) begin
      dat_rsp_l3_pvld <= 1'h0;
    end else begin
      dat_rsp_l3_pvld <= dat_rsp_l2_pvld;
    end
    if (_T_337) begin
      dat_rsp_l1_pvld <= 1'h0;
    end else begin
      dat_rsp_l1_pvld <= dat_rsp_l0_pvld;
    end
    if (_T_337) begin
      dat_rsp_l0_pvld <= 1'h0;
    end else begin
      dat_rsp_l0_pvld <= dat_rsp_pipe_pvld;
    end
    if (_T_337) begin
      _T_1617 <= 27'h0;
    end else begin
      if (dat_rsp_l2_pvld) begin
        _T_1617 <= _T_1614;
      end
    end
    if (_T_337) begin
      _T_1611 <= 27'h0;
    end else begin
      if (dat_rsp_l0_pvld) begin
        _T_1611 <= _T_1608;
      end
    end
    if (_T_337) begin
      _T_1608 <= 27'h0;
    end else begin
      if (dat_rsp_pipe_pvld) begin
        _T_1608 <= _T_1626;
      end
    end
    if (_T_337) begin
      _T_773 <= 1'h0;
    end else begin
      _T_773 <= dat_rls;
    end
    if (_T_337) begin
      _T_776 <= 14'h0;
    end else begin
      if (dat_rls) begin
        if (sub_rls) begin
          _T_776 <= rls_slices;
        end else begin
          _T_776 <= last_slices;
        end
      end
    end
    if (_T_337) begin
      _T_779 <= 15'h0;
    end else begin
      if (dat_rls) begin
        if (sub_rls) begin
          _T_779 <= rls_entries;
        end else begin
          _T_779 <= last_entries;
        end
      end
    end
    if (_T_337) begin
      _T_784 <= 1'h0;
    end else begin
      _T_784 <= sg2dl_pvld;
    end
    if (_T_337) begin
      _T_787 <= 1'h0;
    end else begin
      _T_787 <= _T_784;
    end
    if (_T_337) begin
      _T_790 <= 1'h0;
    end else begin
      _T_790 <= _T_787;
    end
    if (_T_337) begin
      _T_793 <= 1'h0;
    end else begin
      _T_793 <= _T_790;
    end
    if (_T_337) begin
      dl_in_pvld <= 1'h0;
    end else begin
      dl_in_pvld <= _T_793;
    end
    if (_T_337) begin
      _T_817 <= 1'h0;
    end else begin
      _T_817 <= dl_in_pvld;
    end
    if (_T_337) begin
      _T_820 <= 1'h0;
    end else begin
      _T_820 <= _T_817;
    end
    if (_T_337) begin
      _T_823 <= 1'h0;
    end else begin
      _T_823 <= _T_820;
    end
    if (_T_337) begin
      _T_826 <= 1'h0;
    end else begin
      _T_826 <= _T_823;
    end
    if (_T_337) begin
      _T_831 <= 31'h0;
    end else begin
      if (dl_in_pvld) begin
        _T_831 <= _T_828;
      end
    end
    if (_T_337) begin
      _T_834 <= 31'h0;
    end else begin
      if (_T_817) begin
        _T_834 <= _T_831;
      end
    end
    if (_T_337) begin
      _T_837 <= 31'h0;
    end else begin
      if (_T_820) begin
        _T_837 <= _T_834;
      end
    end
    if (_T_337) begin
      _T_840 <= 31'h0;
    end else begin
      if (_T_823) begin
        _T_840 <= _T_837;
      end
    end
    if (_T_337) begin
      batch_cnt <= 6'h0;
    end else begin
      batch_cnt <= _T_877;
    end
    if (_T_337) begin
      sub_h_cnt <= 2'h0;
    end else begin
      sub_h_cnt <= _GEN_65[1:0];
    end
    if (_T_337) begin
      stripe_cnt <= 7'h0;
    end else begin
      stripe_cnt <= _GEN_66[6:0];
    end
    if (_T_337) begin
      dat_exec_valid_d1 <= 1'h0;
    end else begin
      if (dl_pvld) begin
        dat_exec_valid_d1 <= 1'h1;
      end else begin
        if (_T_930) begin
          dat_exec_valid_d1 <= 1'h0;
        end
      end
    end
    if (_T_337) begin
      dat_pipe_local_valid <= 1'h0;
    end else begin
      if (_T_914) begin
        dat_pipe_local_valid <= 1'h0;
      end else begin
        if (dl_pvld) begin
          dat_pipe_local_valid <= 1'h1;
        end
      end
    end
    if (_T_337) begin
      dat_pipe_valid_d1 <= 1'h0;
    end else begin
      dat_pipe_valid_d1 <= dat_pipe_valid;
    end
    if (_T_337) begin
      dat_req_bytes_d1 <= 8'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_bytes_d1 <= dat_req_bytes;
      end
    end
    if (_T_337) begin
      dataout_w_cnt <= 13'h0;
    end else begin
      if (dataout_w_cnt_reg_en) begin
        if (layer_st) begin
          dataout_w_cnt <= {{9'd0}, dataout_w_init};
        end else begin
          if (_T_946) begin
            dataout_w_cnt <= dataout_w_ori;
          end else begin
            if (is_w_end) begin
              dataout_w_cnt <= {{9'd0}, dataout_w_init};
            end else begin
              dataout_w_cnt <= dataout_w_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      dataout_w_ori <= 13'h0;
    end else begin
      if (dataout_w_ori_reg_en) begin
        if (layer_st) begin
          dataout_w_ori <= {{9'd0}, dataout_w_init};
        end else begin
          if (!(_T_946)) begin
            if (is_w_end) begin
              dataout_w_ori <= {{9'd0}, dataout_w_init};
            end else begin
              dataout_w_ori <= dataout_w_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      datain_c_cnt <= 11'h0;
    end else begin
      if (datain_c_cnt_reg_en) begin
        if (layer_st) begin
          datain_c_cnt <= 11'h0;
        end else begin
          if (dl_channel_end) begin
            datain_c_cnt <= 11'h0;
          end else begin
            datain_c_cnt <= _T_961;
          end
        end
      end
    end
    if (_T_337) begin
      datain_w_cnt <= 14'h0;
    end else begin
      if (datain_w_cnt_reg_en) begin
        if (layer_st) begin
          if (is_img) begin
            datain_w_cnt <= 14'h0;
          end else begin
            datain_w_cnt <= _T_984;
          end
        end else begin
          if (_T_946) begin
            datain_w_cnt <= datain_w_ori;
          end else begin
            if (is_w_end) begin
              if (is_img) begin
                datain_w_cnt <= 14'h0;
              end else begin
                datain_w_cnt <= _T_984;
              end
            end else begin
              datain_w_cnt <= datain_w_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      datain_w_ori <= 14'h0;
    end else begin
      if (datain_w_ori_reg_en) begin
        if (layer_st) begin
          if (is_img) begin
            datain_w_ori <= 14'h0;
          end else begin
            datain_w_ori <= _T_984;
          end
        end else begin
          if (!(_T_946)) begin
            if (is_w_end) begin
              if (is_img) begin
                datain_w_ori <= 14'h0;
              end else begin
                datain_w_ori <= _T_984;
              end
            end else begin
              datain_w_ori <= datain_w_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      pixel_w_cnt <= 16'h0;
    end else begin
      if (datain_w_cnt_reg_en) begin
        pixel_w_cnt <= pixel_w_cnt_w;
      end
    end
    if (_T_337) begin
      pixel_w_ori <= 16'h0;
    end else begin
      if (datain_w_ori_reg_en) begin
        pixel_w_ori <= pixel_w_cnt_w;
      end
    end
    if (_T_337) begin
      pixel_w_ch_ori <= 16'h0;
    end else begin
      if (pixel_ch_ori_reg_en) begin
        pixel_w_ch_ori <= pixel_w_cnt_w;
      end
    end
    if (_T_337) begin
      channel_op_cnt <= 13'h2;
    end else begin
      channel_op_cnt <= _T_1016[12:0];
    end
    if (_T_337) begin
      pixel_force_clr_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        pixel_force_clr_d1 <= pixel_force_clr;
      end
    end
    if (_T_337) begin
      pixel_force_fetch_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        if (_T_1062) begin
          pixel_force_fetch_d1 <= 1'h1;
        end else begin
          if (pixel_force_clr_d1) begin
            pixel_force_fetch_d1 <= 1'h0;
          end
        end
      end
    end
    if (_T_337) begin
      datain_h_cnt <= 14'h0;
    end else begin
      if (datain_h_cnt_reg_en) begin
        if (_T_1078) begin
          datain_h_cnt <= datain_h_cnt_st;
        end else begin
          if (_T_946) begin
            datain_h_cnt <= datain_h_ori;
          end else begin
            if (is_w_end) begin
              datain_h_cnt <= datain_h_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      datain_h_ori <= 14'h0;
    end else begin
      if (dataout_w_ori_reg_en) begin
        if (_T_1078) begin
          datain_h_ori <= datain_h_cnt_st;
        end else begin
          if (!(_T_946)) begin
            if (is_w_end) begin
              datain_h_ori <= datain_h_cnt_inc;
            end else begin
              datain_h_ori <= datain_h_cnt;
            end
          end
        end
      end
    end
    if (_T_337) begin
      dat_req_valid_d1 <= 1'h0;
    end else begin
      dat_req_valid_d1 <= dat_req_valid;
    end
    if (_T_337) begin
      dat_req_sub_w_d1 <= 2'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_sub_w_d1 <= dat_req_sub_w_w;
      end
    end
    if (_T_337) begin
      dat_req_sub_h_d1 <= 2'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_sub_h_d1 <= sub_h_cnt;
      end
    end
    if (_T_337) begin
      dat_req_sub_c_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        if (_T_1115) begin
          dat_req_sub_c_d1 <= _T_1116;
        end else begin
          dat_req_sub_c_d1 <= dl_block_end;
        end
      end
    end
    if (_T_337) begin
      dat_req_ch_end_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_ch_end_d1 <= is_last_channel;
      end
    end
    if (_T_337) begin
      dat_req_dummy_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        if (dl_pvld) begin
          dat_req_dummy_d1 <= 1'h1;
        end else begin
          if (_T_930) begin
            dat_req_dummy_d1 <= 1'h0;
          end else begin
            dat_req_dummy_d1 <= dat_exec_valid_d1;
          end
        end
      end
    end
    if (_T_337) begin
      dat_req_cur_sub_h_d1 <= 2'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_cur_sub_h_d1 <= dl_cur_sub_h;
      end
    end
    if (_T_337) begin
      dat_req_sub_w_st_d1 <= 1'h0;
    end else begin
      if (dat_req_sub_w_st_en) begin
        dat_req_sub_w_st_d1 <= dl_pvld;
      end
    end
    if (_T_337) begin
      dat_req_flag_d1 <= 9'h0;
    end else begin
      dat_req_flag_d1 <= _GEN_84[8:0];
    end
    if (_T_337) begin
      dat_req_rls_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_rls_d1 <= _T_1143;
      end
    end
    if (_T_337) begin
      c_bias <= 13'h0;
    end else begin
      if (datain_c_cnt_reg_en) begin
        if (layer_st) begin
          c_bias <= 13'h0;
        end else begin
          if (_T_1163) begin
            c_bias <= 13'h0;
          end else begin
            c_bias <= _T_1166;
          end
        end
      end
    end
    if (_T_337) begin
      c_bias_d1 <= 13'h0;
    end else begin
      if (c_bias_d1_reg_en) begin
        c_bias_d1 <= c_bias;
      end
    end
    if (_T_337) begin
      h_bias_0_d1 <= 13'h0;
    end else begin
      if (_T_1196) begin
        h_bias_0_d1 <= h_bias_0_w;
      end
    end
    if (_T_337) begin
      h_bias_1_d1 <= 13'h0;
    end else begin
      if (_T_1196) begin
        h_bias_1_d1 <= h_bias_1_w;
      end
    end
    if (_T_337) begin
      h_bias_2_d1 <= 13'h0;
    end else begin
      if (_T_1196) begin
        h_bias_2_d1 <= h_bias_2_w;
      end
    end
    if (_T_337) begin
      h_bias_3_d1 <= 13'h0;
    end else begin
      if (_T_1197) begin
        h_bias_3_d1 <= h_bias_3_w;
      end
    end
    if (_T_337) begin
      w_bias_d1 <= 13'h0;
    end else begin
      w_bias_d1 <= _GEN_95[12:0];
    end
    if (_T_337) begin
      dat_req_sub_h_addr_0 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_0 <= _GEN_96[12:0];
    end
    if (_T_337) begin
      dat_req_sub_h_addr_1 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_1 <= _GEN_97[12:0];
    end
    if (_T_337) begin
      dat_req_sub_h_addr_2 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_2 <= _GEN_98[12:0];
    end
    if (_T_337) begin
      sc2buf_dat_rd_en_out <= 1'h0;
    end else begin
      sc2buf_dat_rd_en_out <= sc2buf_dat_rd_en_w;
    end
    if (_T_337) begin
      sc2buf_dat_rd_addr_out <= 18'h1fff;
    end else begin
      if (_T_1369) begin
        if (_T_1307) begin
          sc2buf_dat_rd_addr_out <= 18'h1fff;
        end else begin
          if (is_dat_req_addr_wrap) begin
            sc2buf_dat_rd_addr_out <= dat_req_addr_wrap;
          end else begin
            sc2buf_dat_rd_addr_out <= {{5'd0}, _T_1313};
          end
        end
      end
    end
    if (_T_337) begin
      dat_req_pipe_pvld <= 1'h0;
    end else begin
      dat_req_pipe_pvld <= dat_pipe_valid_d1;
    end
    if (_T_337) begin
      dat_req_pipe_sub_w <= 2'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_w <= dat_req_sub_w_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_sub_h <= 2'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_h <= dat_req_sub_h_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_sub_c <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_c <= dat_req_sub_c_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_ch_end <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_ch_end <= dat_req_ch_end_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_bytes <= 8'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_bytes <= dat_req_bytes_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_dummy <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_dummy <= dat_req_dummy_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_cur_sub_h <= 2'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_cur_sub_h <= dat_req_cur_sub_h_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_sub_w_st <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_w_st <= dat_req_sub_w_st_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_rls <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_rls <= dat_req_rls_d1;
      end
    end
    if (_T_337) begin
      dat_req_pipe_flag <= 9'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_flag <= dat_req_flag_d1;
      end else begin
        dat_req_pipe_flag <= {{8'd0}, dat_exec_valid_d1};
      end
    end
    if (_T_337) begin
      _T_1389 <= 1'h0;
    end else begin
      _T_1389 <= dat_req_pipe_pvld;
    end
    if (_T_337) begin
      _T_1392 <= 1'h0;
    end else begin
      _T_1392 <= _T_1389;
    end
    if (_T_337) begin
      _T_1395 <= 1'h0;
    end else begin
      _T_1395 <= _T_1392;
    end
    if (_T_337) begin
      _T_1398 <= 1'h0;
    end else begin
      _T_1398 <= _T_1395;
    end
    if (_T_337) begin
      _T_1401 <= 1'h0;
    end else begin
      _T_1401 <= _T_1398;
    end
    if (_T_337) begin
      dat_rsp_pipe_pvld <= 1'h0;
    end else begin
      dat_rsp_pipe_pvld <= _T_1401;
    end
    if (_T_337) begin
      _T_1408 <= 29'h0;
    end else begin
      if (dat_req_pipe_pvld) begin
        _T_1408 <= dat_req_pipe_pd;
      end
    end
    if (_T_337) begin
      _T_1411 <= 29'h0;
    end else begin
      if (_T_1389) begin
        _T_1411 <= _T_1408;
      end
    end
    if (_T_337) begin
      _T_1414 <= 29'h0;
    end else begin
      if (_T_1392) begin
        _T_1414 <= _T_1411;
      end
    end
    if (_T_337) begin
      _T_1417 <= 29'h0;
    end else begin
      if (_T_1395) begin
        _T_1417 <= _T_1414;
      end
    end
    if (_T_337) begin
      _T_1420 <= 29'h0;
    end else begin
      if (_T_1398) begin
        _T_1420 <= _T_1417;
      end
    end
    if (_T_337) begin
      dat_rsp_pipe_pd <= 29'h0;
    end else begin
      if (_T_1401) begin
        dat_rsp_pipe_pd <= _T_1420;
      end
    end
    if (_T_337) begin
      dat_l0c0_dummy <= 1'h1;
    end else begin
      if (sc2buf_dat_rd_valid) begin
        dat_l0c0_dummy <= 1'h0;
      end
    end
    if (_T_337) begin
      dat_l0c1_dummy <= 1'h1;
    end else begin
      if (dat_l0c1_en) begin
        dat_l0c1_dummy <= 1'h0;
      end else begin
        if (sc2buf_dat_rd_valid) begin
          dat_l0c1_dummy <= dat_l0c0_dummy;
        end
      end
    end
    if (sc2buf_dat_rd_valid) begin
      dat_l0c0 <= sc2buf_dat_rd_data;
    end
    if (dat_l0c1_en) begin
      dat_l0c1 <= dat_l0c0;
    end
    if (_T_337) begin
      rsp_sft_cnt_l0 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l0_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l0 <= 8'h40;
        end else begin
          if (_T_1691) begin
            rsp_sft_cnt_l0 <= rsp_sft_cnt_l0_ori;
          end else begin
            if (_T_1692) begin
              rsp_sft_cnt_l0 <= 8'h40;
            end else begin
              rsp_sft_cnt_l0 <= rsp_sft_cnt_l0_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l1 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l1_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l1 <= 8'h40;
        end else begin
          if (_T_1701) begin
            rsp_sft_cnt_l1 <= rsp_sft_cnt_l1_ori;
          end else begin
            if (_T_1702) begin
              rsp_sft_cnt_l1 <= 8'h40;
            end else begin
              rsp_sft_cnt_l1 <= rsp_sft_cnt_l1_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l2 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l2_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l2 <= 8'h40;
        end else begin
          if (_T_1711) begin
            rsp_sft_cnt_l2 <= rsp_sft_cnt_l2_ori;
          end else begin
            if (_T_1712) begin
              rsp_sft_cnt_l2 <= 8'h40;
            end else begin
              rsp_sft_cnt_l2 <= rsp_sft_cnt_l2_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l3 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l3_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l3 <= 8'h40;
        end else begin
          if (_T_1721) begin
            rsp_sft_cnt_l3 <= rsp_sft_cnt_l3_ori;
          end else begin
            if (_T_1722) begin
              rsp_sft_cnt_l3 <= 8'h40;
            end else begin
              rsp_sft_cnt_l3 <= rsp_sft_cnt_l3_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l0_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l0_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l0_ori <= 8'h40;
        end else begin
          if (!(_T_1691)) begin
            if (_T_1692) begin
              rsp_sft_cnt_l0_ori <= 8'h40;
            end else begin
              rsp_sft_cnt_l0_ori <= rsp_sft_cnt_l0_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l1_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l1_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l1_ori <= 8'h40;
        end else begin
          if (!(_T_1701)) begin
            if (_T_1702) begin
              rsp_sft_cnt_l1_ori <= 8'h40;
            end else begin
              rsp_sft_cnt_l1_ori <= rsp_sft_cnt_l1_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l2_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l2_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l2_ori <= 8'h40;
        end else begin
          if (!(_T_1711)) begin
            if (_T_1712) begin
              rsp_sft_cnt_l2_ori <= 8'h40;
            end else begin
              rsp_sft_cnt_l2_ori <= rsp_sft_cnt_l2_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      rsp_sft_cnt_l3_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l3_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l3_ori <= 8'h40;
        end else begin
          if (!(_T_1721)) begin
            if (_T_1722) begin
              rsp_sft_cnt_l3_ori <= 8'h40;
            end else begin
              rsp_sft_cnt_l3_ori <= rsp_sft_cnt_l3_inc;
            end
          end
        end
      end
    end
    if (_T_337) begin
      dat_rsp_l2_pvld <= 1'h0;
    end else begin
      dat_rsp_l2_pvld <= dat_rsp_l1_pvld;
    end
    if (_T_337) begin
      _T_1614 <= 27'h0;
    end else begin
      if (dat_rsp_l1_pvld) begin
        _T_1614 <= _T_1611;
      end
    end
    dat_rsp_l0_sft_d1 <= _GEN_149[255:0];
    dat_rsp_l0_sft_d2 <= _GEN_150[127:0];
    if (dat_rsp_sft_d3_en) begin
      dat_rsp_l0_sft_d3 <= dat_rsp_l0_sft_d2;
    end
    dat_rsp_l1_sft_d2 <= _GEN_151[127:0];
    if (dat_rsp_sft_d3_en) begin
      dat_rsp_l1_sft_d3 <= dat_rsp_l1_sft_d2;
    end
    dat_rsp_l2_sft_d3 <= _GEN_154[127:0];
    if (_T_337) begin
      dat_out_pvld <= 1'h0;
    end else begin
      dat_out_pvld <= dat_rsp_pvld;
    end
    if (_T_337) begin
      dat_out_flag <= 9'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_flag <= dat_rsp_flag;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_0 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_0 <= dat_rsp_mask_w_0;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_1 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_1 <= dat_rsp_mask_w_1;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_2 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_2 <= dat_rsp_mask_w_2;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_3 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_3 <= dat_rsp_mask_w_3;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_4 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_4 <= dat_rsp_mask_w_4;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_5 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_5 <= dat_rsp_mask_w_5;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_6 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_6 <= dat_rsp_mask_w_6;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_7 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_7 <= dat_rsp_mask_w_7;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_8 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_8 <= dat_rsp_mask_w_8;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_9 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_9 <= dat_rsp_mask_w_9;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_10 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_10 <= dat_rsp_mask_w_10;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_11 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_11 <= dat_rsp_mask_w_11;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_12 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_12 <= dat_rsp_mask_w_12;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_13 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_13 <= dat_rsp_mask_w_13;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_14 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_14 <= dat_rsp_mask_w_14;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_15 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_15 <= dat_rsp_mask_w_15;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_16 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_16 <= dat_rsp_mask_w_16;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_17 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_17 <= dat_rsp_mask_w_17;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_18 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_18 <= dat_rsp_mask_w_18;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_19 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_19 <= dat_rsp_mask_w_19;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_20 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_20 <= dat_rsp_mask_w_20;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_21 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_21 <= dat_rsp_mask_w_21;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_22 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_22 <= dat_rsp_mask_w_22;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_23 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_23 <= dat_rsp_mask_w_23;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_24 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_24 <= dat_rsp_mask_w_24;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_25 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_25 <= dat_rsp_mask_w_25;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_26 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_26 <= dat_rsp_mask_w_26;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_27 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_27 <= dat_rsp_mask_w_27;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_28 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_28 <= dat_rsp_mask_w_28;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_29 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_29 <= dat_rsp_mask_w_29;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_30 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_30 <= dat_rsp_mask_w_30;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_31 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_31 <= dat_rsp_mask_w_31;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_32 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_32 <= dat_rsp_mask_w_32;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_33 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_33 <= dat_rsp_mask_w_33;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_34 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_34 <= dat_rsp_mask_w_34;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_35 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_35 <= dat_rsp_mask_w_35;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_36 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_36 <= dat_rsp_mask_w_36;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_37 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_37 <= dat_rsp_mask_w_37;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_38 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_38 <= dat_rsp_mask_w_38;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_39 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_39 <= dat_rsp_mask_w_39;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_40 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_40 <= dat_rsp_mask_w_40;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_41 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_41 <= dat_rsp_mask_w_41;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_42 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_42 <= dat_rsp_mask_w_42;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_43 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_43 <= dat_rsp_mask_w_43;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_44 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_44 <= dat_rsp_mask_w_44;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_45 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_45 <= dat_rsp_mask_w_45;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_46 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_46 <= dat_rsp_mask_w_46;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_47 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_47 <= dat_rsp_mask_w_47;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_48 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_48 <= dat_rsp_mask_w_48;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_49 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_49 <= dat_rsp_mask_w_49;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_50 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_50 <= dat_rsp_mask_w_50;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_51 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_51 <= dat_rsp_mask_w_51;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_52 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_52 <= dat_rsp_mask_w_52;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_53 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_53 <= dat_rsp_mask_w_53;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_54 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_54 <= dat_rsp_mask_w_54;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_55 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_55 <= dat_rsp_mask_w_55;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_56 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_56 <= dat_rsp_mask_w_56;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_57 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_57 <= dat_rsp_mask_w_57;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_58 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_58 <= dat_rsp_mask_w_58;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_59 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_59 <= dat_rsp_mask_w_59;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_60 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_60 <= dat_rsp_mask_w_60;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_61 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_61 <= dat_rsp_mask_w_61;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_62 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_62 <= dat_rsp_mask_w_62;
      end
    end
    if (_T_337) begin
      dat_out_bypass_mask_63 <= 1'h0;
    end else begin
      if (dat_rsp_pvld) begin
        dat_out_bypass_mask_63 <= dat_rsp_mask_w_63;
      end
    end
    if (_T_3247) begin
      if (_T_2186) begin
        dat_out_bypass_data_0 <= dat_rsp_img_0;
      end else begin
        dat_out_bypass_data_0 <= dat_rsp_conv_0;
      end
    end
    if (_T_3248) begin
      if (_T_2186) begin
        dat_out_bypass_data_1 <= dat_rsp_img_1;
      end else begin
        dat_out_bypass_data_1 <= dat_rsp_conv_1;
      end
    end
    if (_T_3249) begin
      if (_T_2186) begin
        dat_out_bypass_data_2 <= dat_rsp_img_2;
      end else begin
        dat_out_bypass_data_2 <= dat_rsp_conv_2;
      end
    end
    if (_T_3250) begin
      if (_T_2186) begin
        dat_out_bypass_data_3 <= dat_rsp_img_3;
      end else begin
        dat_out_bypass_data_3 <= dat_rsp_conv_3;
      end
    end
    if (_T_3251) begin
      if (_T_2186) begin
        dat_out_bypass_data_4 <= dat_rsp_img_4;
      end else begin
        dat_out_bypass_data_4 <= dat_rsp_conv_4;
      end
    end
    if (_T_3252) begin
      if (_T_2186) begin
        dat_out_bypass_data_5 <= dat_rsp_img_5;
      end else begin
        dat_out_bypass_data_5 <= dat_rsp_conv_5;
      end
    end
    if (_T_3253) begin
      if (_T_2186) begin
        dat_out_bypass_data_6 <= dat_rsp_img_6;
      end else begin
        dat_out_bypass_data_6 <= dat_rsp_conv_6;
      end
    end
    if (_T_3254) begin
      if (_T_2186) begin
        dat_out_bypass_data_7 <= dat_rsp_img_7;
      end else begin
        dat_out_bypass_data_7 <= dat_rsp_conv_7;
      end
    end
    if (_T_3255) begin
      if (_T_2186) begin
        dat_out_bypass_data_8 <= dat_rsp_img_8;
      end else begin
        dat_out_bypass_data_8 <= dat_rsp_conv_8;
      end
    end
    if (_T_3256) begin
      if (_T_2186) begin
        dat_out_bypass_data_9 <= dat_rsp_img_9;
      end else begin
        dat_out_bypass_data_9 <= dat_rsp_conv_9;
      end
    end
    if (_T_3257) begin
      if (_T_2186) begin
        dat_out_bypass_data_10 <= dat_rsp_img_10;
      end else begin
        dat_out_bypass_data_10 <= dat_rsp_conv_10;
      end
    end
    if (_T_3258) begin
      if (_T_2186) begin
        dat_out_bypass_data_11 <= dat_rsp_img_11;
      end else begin
        dat_out_bypass_data_11 <= dat_rsp_conv_11;
      end
    end
    if (_T_3259) begin
      if (_T_2186) begin
        dat_out_bypass_data_12 <= dat_rsp_img_12;
      end else begin
        dat_out_bypass_data_12 <= dat_rsp_conv_12;
      end
    end
    if (_T_3260) begin
      if (_T_2186) begin
        dat_out_bypass_data_13 <= dat_rsp_img_13;
      end else begin
        dat_out_bypass_data_13 <= dat_rsp_conv_13;
      end
    end
    if (_T_3261) begin
      if (_T_2186) begin
        dat_out_bypass_data_14 <= dat_rsp_img_14;
      end else begin
        dat_out_bypass_data_14 <= dat_rsp_conv_14;
      end
    end
    if (_T_3262) begin
      if (_T_2186) begin
        dat_out_bypass_data_15 <= dat_rsp_img_15;
      end else begin
        dat_out_bypass_data_15 <= dat_rsp_conv_15;
      end
    end
    if (_T_3263) begin
      if (_T_2186) begin
        dat_out_bypass_data_16 <= dat_rsp_img_16;
      end else begin
        dat_out_bypass_data_16 <= dat_rsp_conv_16;
      end
    end
    if (_T_3264) begin
      if (_T_2186) begin
        dat_out_bypass_data_17 <= dat_rsp_img_17;
      end else begin
        dat_out_bypass_data_17 <= dat_rsp_conv_17;
      end
    end
    if (_T_3265) begin
      if (_T_2186) begin
        dat_out_bypass_data_18 <= dat_rsp_img_18;
      end else begin
        dat_out_bypass_data_18 <= dat_rsp_conv_18;
      end
    end
    if (_T_3266) begin
      if (_T_2186) begin
        dat_out_bypass_data_19 <= dat_rsp_img_19;
      end else begin
        dat_out_bypass_data_19 <= dat_rsp_conv_19;
      end
    end
    if (_T_3267) begin
      if (_T_2186) begin
        dat_out_bypass_data_20 <= dat_rsp_img_20;
      end else begin
        dat_out_bypass_data_20 <= dat_rsp_conv_20;
      end
    end
    if (_T_3268) begin
      if (_T_2186) begin
        dat_out_bypass_data_21 <= dat_rsp_img_21;
      end else begin
        dat_out_bypass_data_21 <= dat_rsp_conv_21;
      end
    end
    if (_T_3269) begin
      if (_T_2186) begin
        dat_out_bypass_data_22 <= dat_rsp_img_22;
      end else begin
        dat_out_bypass_data_22 <= dat_rsp_conv_22;
      end
    end
    if (_T_3270) begin
      if (_T_2186) begin
        dat_out_bypass_data_23 <= dat_rsp_img_23;
      end else begin
        dat_out_bypass_data_23 <= dat_rsp_conv_23;
      end
    end
    if (_T_3271) begin
      if (_T_2186) begin
        dat_out_bypass_data_24 <= dat_rsp_img_24;
      end else begin
        dat_out_bypass_data_24 <= dat_rsp_conv_24;
      end
    end
    if (_T_3272) begin
      if (_T_2186) begin
        dat_out_bypass_data_25 <= dat_rsp_img_25;
      end else begin
        dat_out_bypass_data_25 <= dat_rsp_conv_25;
      end
    end
    if (_T_3273) begin
      if (_T_2186) begin
        dat_out_bypass_data_26 <= dat_rsp_img_26;
      end else begin
        dat_out_bypass_data_26 <= dat_rsp_conv_26;
      end
    end
    if (_T_3274) begin
      if (_T_2186) begin
        dat_out_bypass_data_27 <= dat_rsp_img_27;
      end else begin
        dat_out_bypass_data_27 <= dat_rsp_conv_27;
      end
    end
    if (_T_3275) begin
      if (_T_2186) begin
        dat_out_bypass_data_28 <= dat_rsp_img_28;
      end else begin
        dat_out_bypass_data_28 <= dat_rsp_conv_28;
      end
    end
    if (_T_3276) begin
      if (_T_2186) begin
        dat_out_bypass_data_29 <= dat_rsp_img_29;
      end else begin
        dat_out_bypass_data_29 <= dat_rsp_conv_29;
      end
    end
    if (_T_3277) begin
      if (_T_2186) begin
        dat_out_bypass_data_30 <= dat_rsp_img_30;
      end else begin
        dat_out_bypass_data_30 <= dat_rsp_conv_30;
      end
    end
    if (_T_3278) begin
      if (_T_2186) begin
        dat_out_bypass_data_31 <= dat_rsp_img_31;
      end else begin
        dat_out_bypass_data_31 <= dat_rsp_conv_31;
      end
    end
    if (_T_3279) begin
      if (_T_2186) begin
        dat_out_bypass_data_32 <= dat_rsp_img_32;
      end else begin
        dat_out_bypass_data_32 <= dat_rsp_conv_32;
      end
    end
    if (_T_3280) begin
      if (_T_2186) begin
        dat_out_bypass_data_33 <= dat_rsp_img_33;
      end else begin
        dat_out_bypass_data_33 <= dat_rsp_conv_33;
      end
    end
    if (_T_3281) begin
      if (_T_2186) begin
        dat_out_bypass_data_34 <= dat_rsp_img_34;
      end else begin
        dat_out_bypass_data_34 <= dat_rsp_conv_34;
      end
    end
    if (_T_3282) begin
      if (_T_2186) begin
        dat_out_bypass_data_35 <= dat_rsp_img_35;
      end else begin
        dat_out_bypass_data_35 <= dat_rsp_conv_35;
      end
    end
    if (_T_3283) begin
      if (_T_2186) begin
        dat_out_bypass_data_36 <= dat_rsp_img_36;
      end else begin
        dat_out_bypass_data_36 <= dat_rsp_conv_36;
      end
    end
    if (_T_3284) begin
      if (_T_2186) begin
        dat_out_bypass_data_37 <= dat_rsp_img_37;
      end else begin
        dat_out_bypass_data_37 <= dat_rsp_conv_37;
      end
    end
    if (_T_3285) begin
      if (_T_2186) begin
        dat_out_bypass_data_38 <= dat_rsp_img_38;
      end else begin
        dat_out_bypass_data_38 <= dat_rsp_conv_38;
      end
    end
    if (_T_3286) begin
      if (_T_2186) begin
        dat_out_bypass_data_39 <= dat_rsp_img_39;
      end else begin
        dat_out_bypass_data_39 <= dat_rsp_conv_39;
      end
    end
    if (_T_3287) begin
      if (_T_2186) begin
        dat_out_bypass_data_40 <= dat_rsp_img_40;
      end else begin
        dat_out_bypass_data_40 <= dat_rsp_conv_40;
      end
    end
    if (_T_3288) begin
      if (_T_2186) begin
        dat_out_bypass_data_41 <= dat_rsp_img_41;
      end else begin
        dat_out_bypass_data_41 <= dat_rsp_conv_41;
      end
    end
    if (_T_3289) begin
      if (_T_2186) begin
        dat_out_bypass_data_42 <= dat_rsp_img_42;
      end else begin
        dat_out_bypass_data_42 <= dat_rsp_conv_42;
      end
    end
    if (_T_3290) begin
      if (_T_2186) begin
        dat_out_bypass_data_43 <= dat_rsp_img_43;
      end else begin
        dat_out_bypass_data_43 <= dat_rsp_conv_43;
      end
    end
    if (_T_3291) begin
      if (_T_2186) begin
        dat_out_bypass_data_44 <= dat_rsp_img_44;
      end else begin
        dat_out_bypass_data_44 <= dat_rsp_conv_44;
      end
    end
    if (_T_3292) begin
      if (_T_2186) begin
        dat_out_bypass_data_45 <= dat_rsp_img_45;
      end else begin
        dat_out_bypass_data_45 <= dat_rsp_conv_45;
      end
    end
    if (_T_3293) begin
      if (_T_2186) begin
        dat_out_bypass_data_46 <= dat_rsp_img_46;
      end else begin
        dat_out_bypass_data_46 <= dat_rsp_conv_46;
      end
    end
    if (_T_3294) begin
      if (_T_2186) begin
        dat_out_bypass_data_47 <= dat_rsp_img_47;
      end else begin
        dat_out_bypass_data_47 <= dat_rsp_conv_47;
      end
    end
    if (_T_3295) begin
      if (_T_2186) begin
        dat_out_bypass_data_48 <= dat_rsp_img_48;
      end else begin
        dat_out_bypass_data_48 <= dat_rsp_conv_48;
      end
    end
    if (_T_3296) begin
      if (_T_2186) begin
        dat_out_bypass_data_49 <= dat_rsp_img_49;
      end else begin
        dat_out_bypass_data_49 <= dat_rsp_conv_49;
      end
    end
    if (_T_3297) begin
      if (_T_2186) begin
        dat_out_bypass_data_50 <= dat_rsp_img_50;
      end else begin
        dat_out_bypass_data_50 <= dat_rsp_conv_50;
      end
    end
    if (_T_3298) begin
      if (_T_2186) begin
        dat_out_bypass_data_51 <= dat_rsp_img_51;
      end else begin
        dat_out_bypass_data_51 <= dat_rsp_conv_51;
      end
    end
    if (_T_3299) begin
      if (_T_2186) begin
        dat_out_bypass_data_52 <= dat_rsp_img_52;
      end else begin
        dat_out_bypass_data_52 <= dat_rsp_conv_52;
      end
    end
    if (_T_3300) begin
      if (_T_2186) begin
        dat_out_bypass_data_53 <= dat_rsp_img_53;
      end else begin
        dat_out_bypass_data_53 <= dat_rsp_conv_53;
      end
    end
    if (_T_3301) begin
      if (_T_2186) begin
        dat_out_bypass_data_54 <= dat_rsp_img_54;
      end else begin
        dat_out_bypass_data_54 <= dat_rsp_conv_54;
      end
    end
    if (_T_3302) begin
      if (_T_2186) begin
        dat_out_bypass_data_55 <= dat_rsp_img_55;
      end else begin
        dat_out_bypass_data_55 <= dat_rsp_conv_55;
      end
    end
    if (_T_3303) begin
      if (_T_2186) begin
        dat_out_bypass_data_56 <= dat_rsp_img_56;
      end else begin
        dat_out_bypass_data_56 <= dat_rsp_conv_56;
      end
    end
    if (_T_3304) begin
      if (_T_2186) begin
        dat_out_bypass_data_57 <= dat_rsp_img_57;
      end else begin
        dat_out_bypass_data_57 <= dat_rsp_conv_57;
      end
    end
    if (_T_3305) begin
      if (_T_2186) begin
        dat_out_bypass_data_58 <= dat_rsp_img_58;
      end else begin
        dat_out_bypass_data_58 <= dat_rsp_conv_58;
      end
    end
    if (_T_3306) begin
      if (_T_2186) begin
        dat_out_bypass_data_59 <= dat_rsp_img_59;
      end else begin
        dat_out_bypass_data_59 <= dat_rsp_conv_59;
      end
    end
    if (_T_3307) begin
      if (_T_2186) begin
        dat_out_bypass_data_60 <= dat_rsp_img_60;
      end else begin
        dat_out_bypass_data_60 <= dat_rsp_conv_60;
      end
    end
    if (_T_3308) begin
      if (_T_2186) begin
        dat_out_bypass_data_61 <= dat_rsp_img_61;
      end else begin
        dat_out_bypass_data_61 <= dat_rsp_conv_61;
      end
    end
    if (_T_3309) begin
      if (_T_2186) begin
        dat_out_bypass_data_62 <= dat_rsp_img_62;
      end else begin
        dat_out_bypass_data_62 <= dat_rsp_conv_62;
      end
    end
    if (_T_3310) begin
      if (_T_2186) begin
        dat_out_bypass_data_63 <= dat_rsp_img_63;
      end else begin
        dat_out_bypass_data_63 <= dat_rsp_conv_63;
      end
    end
    if (_T_337) begin
      dl_out_pvld <= 1'h0;
    end else begin
      dl_out_pvld <= dat_out_pvld;
    end
    if (_T_337) begin
      dl_out_mask_0 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_0 <= 1'h0;
        end else begin
          dl_out_mask_0 <= dat_out_bypass_mask_0;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_1 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_1 <= 1'h0;
        end else begin
          dl_out_mask_1 <= dat_out_bypass_mask_1;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_2 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_2 <= 1'h0;
        end else begin
          dl_out_mask_2 <= dat_out_bypass_mask_2;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_3 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_3 <= 1'h0;
        end else begin
          dl_out_mask_3 <= dat_out_bypass_mask_3;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_4 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_4 <= 1'h0;
        end else begin
          dl_out_mask_4 <= dat_out_bypass_mask_4;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_5 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_5 <= 1'h0;
        end else begin
          dl_out_mask_5 <= dat_out_bypass_mask_5;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_6 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_6 <= 1'h0;
        end else begin
          dl_out_mask_6 <= dat_out_bypass_mask_6;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_7 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_7 <= 1'h0;
        end else begin
          dl_out_mask_7 <= dat_out_bypass_mask_7;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_8 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_8 <= 1'h0;
        end else begin
          dl_out_mask_8 <= dat_out_bypass_mask_8;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_9 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_9 <= 1'h0;
        end else begin
          dl_out_mask_9 <= dat_out_bypass_mask_9;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_10 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_10 <= 1'h0;
        end else begin
          dl_out_mask_10 <= dat_out_bypass_mask_10;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_11 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_11 <= 1'h0;
        end else begin
          dl_out_mask_11 <= dat_out_bypass_mask_11;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_12 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_12 <= 1'h0;
        end else begin
          dl_out_mask_12 <= dat_out_bypass_mask_12;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_13 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_13 <= 1'h0;
        end else begin
          dl_out_mask_13 <= dat_out_bypass_mask_13;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_14 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_14 <= 1'h0;
        end else begin
          dl_out_mask_14 <= dat_out_bypass_mask_14;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_15 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_15 <= 1'h0;
        end else begin
          dl_out_mask_15 <= dat_out_bypass_mask_15;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_16 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_16 <= 1'h0;
        end else begin
          dl_out_mask_16 <= dat_out_bypass_mask_16;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_17 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_17 <= 1'h0;
        end else begin
          dl_out_mask_17 <= dat_out_bypass_mask_17;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_18 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_18 <= 1'h0;
        end else begin
          dl_out_mask_18 <= dat_out_bypass_mask_18;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_19 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_19 <= 1'h0;
        end else begin
          dl_out_mask_19 <= dat_out_bypass_mask_19;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_20 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_20 <= 1'h0;
        end else begin
          dl_out_mask_20 <= dat_out_bypass_mask_20;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_21 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_21 <= 1'h0;
        end else begin
          dl_out_mask_21 <= dat_out_bypass_mask_21;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_22 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_22 <= 1'h0;
        end else begin
          dl_out_mask_22 <= dat_out_bypass_mask_22;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_23 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_23 <= 1'h0;
        end else begin
          dl_out_mask_23 <= dat_out_bypass_mask_23;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_24 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_24 <= 1'h0;
        end else begin
          dl_out_mask_24 <= dat_out_bypass_mask_24;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_25 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_25 <= 1'h0;
        end else begin
          dl_out_mask_25 <= dat_out_bypass_mask_25;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_26 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_26 <= 1'h0;
        end else begin
          dl_out_mask_26 <= dat_out_bypass_mask_26;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_27 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_27 <= 1'h0;
        end else begin
          dl_out_mask_27 <= dat_out_bypass_mask_27;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_28 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_28 <= 1'h0;
        end else begin
          dl_out_mask_28 <= dat_out_bypass_mask_28;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_29 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_29 <= 1'h0;
        end else begin
          dl_out_mask_29 <= dat_out_bypass_mask_29;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_30 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_30 <= 1'h0;
        end else begin
          dl_out_mask_30 <= dat_out_bypass_mask_30;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_31 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_31 <= 1'h0;
        end else begin
          dl_out_mask_31 <= dat_out_bypass_mask_31;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_32 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_32 <= 1'h0;
        end else begin
          dl_out_mask_32 <= dat_out_bypass_mask_32;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_33 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_33 <= 1'h0;
        end else begin
          dl_out_mask_33 <= dat_out_bypass_mask_33;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_34 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_34 <= 1'h0;
        end else begin
          dl_out_mask_34 <= dat_out_bypass_mask_34;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_35 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_35 <= 1'h0;
        end else begin
          dl_out_mask_35 <= dat_out_bypass_mask_35;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_36 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_36 <= 1'h0;
        end else begin
          dl_out_mask_36 <= dat_out_bypass_mask_36;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_37 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_37 <= 1'h0;
        end else begin
          dl_out_mask_37 <= dat_out_bypass_mask_37;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_38 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_38 <= 1'h0;
        end else begin
          dl_out_mask_38 <= dat_out_bypass_mask_38;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_39 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_39 <= 1'h0;
        end else begin
          dl_out_mask_39 <= dat_out_bypass_mask_39;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_40 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_40 <= 1'h0;
        end else begin
          dl_out_mask_40 <= dat_out_bypass_mask_40;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_41 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_41 <= 1'h0;
        end else begin
          dl_out_mask_41 <= dat_out_bypass_mask_41;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_42 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_42 <= 1'h0;
        end else begin
          dl_out_mask_42 <= dat_out_bypass_mask_42;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_43 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_43 <= 1'h0;
        end else begin
          dl_out_mask_43 <= dat_out_bypass_mask_43;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_44 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_44 <= 1'h0;
        end else begin
          dl_out_mask_44 <= dat_out_bypass_mask_44;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_45 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_45 <= 1'h0;
        end else begin
          dl_out_mask_45 <= dat_out_bypass_mask_45;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_46 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_46 <= 1'h0;
        end else begin
          dl_out_mask_46 <= dat_out_bypass_mask_46;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_47 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_47 <= 1'h0;
        end else begin
          dl_out_mask_47 <= dat_out_bypass_mask_47;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_48 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_48 <= 1'h0;
        end else begin
          dl_out_mask_48 <= dat_out_bypass_mask_48;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_49 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_49 <= 1'h0;
        end else begin
          dl_out_mask_49 <= dat_out_bypass_mask_49;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_50 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_50 <= 1'h0;
        end else begin
          dl_out_mask_50 <= dat_out_bypass_mask_50;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_51 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_51 <= 1'h0;
        end else begin
          dl_out_mask_51 <= dat_out_bypass_mask_51;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_52 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_52 <= 1'h0;
        end else begin
          dl_out_mask_52 <= dat_out_bypass_mask_52;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_53 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_53 <= 1'h0;
        end else begin
          dl_out_mask_53 <= dat_out_bypass_mask_53;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_54 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_54 <= 1'h0;
        end else begin
          dl_out_mask_54 <= dat_out_bypass_mask_54;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_55 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_55 <= 1'h0;
        end else begin
          dl_out_mask_55 <= dat_out_bypass_mask_55;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_56 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_56 <= 1'h0;
        end else begin
          dl_out_mask_56 <= dat_out_bypass_mask_56;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_57 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_57 <= 1'h0;
        end else begin
          dl_out_mask_57 <= dat_out_bypass_mask_57;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_58 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_58 <= 1'h0;
        end else begin
          dl_out_mask_58 <= dat_out_bypass_mask_58;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_59 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_59 <= 1'h0;
        end else begin
          dl_out_mask_59 <= dat_out_bypass_mask_59;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_60 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_60 <= 1'h0;
        end else begin
          dl_out_mask_60 <= dat_out_bypass_mask_60;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_61 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_61 <= 1'h0;
        end else begin
          dl_out_mask_61 <= dat_out_bypass_mask_61;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_62 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_62 <= 1'h0;
        end else begin
          dl_out_mask_62 <= dat_out_bypass_mask_62;
        end
      end
    end
    if (_T_337) begin
      dl_out_mask_63 <= 1'h0;
    end else begin
      if (_T_4112) begin
        if (_T_3846) begin
          dl_out_mask_63 <= 1'h0;
        end else begin
          dl_out_mask_63 <= dat_out_bypass_mask_63;
        end
      end
    end
    if (_T_337) begin
      dl_out_flag <= 9'h0;
    end else begin
      if (dat_out_pvld) begin
        dl_out_flag <= dat_out_flag;
      end
    end
    if (dat_out_mask_0) begin
      dl_out_data_0 <= dat_out_bypass_data_0;
    end
    if (dat_out_mask_1) begin
      dl_out_data_1 <= dat_out_bypass_data_1;
    end
    if (dat_out_mask_2) begin
      dl_out_data_2 <= dat_out_bypass_data_2;
    end
    if (dat_out_mask_3) begin
      dl_out_data_3 <= dat_out_bypass_data_3;
    end
    if (dat_out_mask_4) begin
      dl_out_data_4 <= dat_out_bypass_data_4;
    end
    if (dat_out_mask_5) begin
      dl_out_data_5 <= dat_out_bypass_data_5;
    end
    if (dat_out_mask_6) begin
      dl_out_data_6 <= dat_out_bypass_data_6;
    end
    if (dat_out_mask_7) begin
      dl_out_data_7 <= dat_out_bypass_data_7;
    end
    if (dat_out_mask_8) begin
      dl_out_data_8 <= dat_out_bypass_data_8;
    end
    if (dat_out_mask_9) begin
      dl_out_data_9 <= dat_out_bypass_data_9;
    end
    if (dat_out_mask_10) begin
      dl_out_data_10 <= dat_out_bypass_data_10;
    end
    if (dat_out_mask_11) begin
      dl_out_data_11 <= dat_out_bypass_data_11;
    end
    if (dat_out_mask_12) begin
      dl_out_data_12 <= dat_out_bypass_data_12;
    end
    if (dat_out_mask_13) begin
      dl_out_data_13 <= dat_out_bypass_data_13;
    end
    if (dat_out_mask_14) begin
      dl_out_data_14 <= dat_out_bypass_data_14;
    end
    if (dat_out_mask_15) begin
      dl_out_data_15 <= dat_out_bypass_data_15;
    end
    if (dat_out_mask_16) begin
      dl_out_data_16 <= dat_out_bypass_data_16;
    end
    if (dat_out_mask_17) begin
      dl_out_data_17 <= dat_out_bypass_data_17;
    end
    if (dat_out_mask_18) begin
      dl_out_data_18 <= dat_out_bypass_data_18;
    end
    if (dat_out_mask_19) begin
      dl_out_data_19 <= dat_out_bypass_data_19;
    end
    if (dat_out_mask_20) begin
      dl_out_data_20 <= dat_out_bypass_data_20;
    end
    if (dat_out_mask_21) begin
      dl_out_data_21 <= dat_out_bypass_data_21;
    end
    if (dat_out_mask_22) begin
      dl_out_data_22 <= dat_out_bypass_data_22;
    end
    if (dat_out_mask_23) begin
      dl_out_data_23 <= dat_out_bypass_data_23;
    end
    if (dat_out_mask_24) begin
      dl_out_data_24 <= dat_out_bypass_data_24;
    end
    if (dat_out_mask_25) begin
      dl_out_data_25 <= dat_out_bypass_data_25;
    end
    if (dat_out_mask_26) begin
      dl_out_data_26 <= dat_out_bypass_data_26;
    end
    if (dat_out_mask_27) begin
      dl_out_data_27 <= dat_out_bypass_data_27;
    end
    if (dat_out_mask_28) begin
      dl_out_data_28 <= dat_out_bypass_data_28;
    end
    if (dat_out_mask_29) begin
      dl_out_data_29 <= dat_out_bypass_data_29;
    end
    if (dat_out_mask_30) begin
      dl_out_data_30 <= dat_out_bypass_data_30;
    end
    if (dat_out_mask_31) begin
      dl_out_data_31 <= dat_out_bypass_data_31;
    end
    if (dat_out_mask_32) begin
      dl_out_data_32 <= dat_out_bypass_data_32;
    end
    if (dat_out_mask_33) begin
      dl_out_data_33 <= dat_out_bypass_data_33;
    end
    if (dat_out_mask_34) begin
      dl_out_data_34 <= dat_out_bypass_data_34;
    end
    if (dat_out_mask_35) begin
      dl_out_data_35 <= dat_out_bypass_data_35;
    end
    if (dat_out_mask_36) begin
      dl_out_data_36 <= dat_out_bypass_data_36;
    end
    if (dat_out_mask_37) begin
      dl_out_data_37 <= dat_out_bypass_data_37;
    end
    if (dat_out_mask_38) begin
      dl_out_data_38 <= dat_out_bypass_data_38;
    end
    if (dat_out_mask_39) begin
      dl_out_data_39 <= dat_out_bypass_data_39;
    end
    if (dat_out_mask_40) begin
      dl_out_data_40 <= dat_out_bypass_data_40;
    end
    if (dat_out_mask_41) begin
      dl_out_data_41 <= dat_out_bypass_data_41;
    end
    if (dat_out_mask_42) begin
      dl_out_data_42 <= dat_out_bypass_data_42;
    end
    if (dat_out_mask_43) begin
      dl_out_data_43 <= dat_out_bypass_data_43;
    end
    if (dat_out_mask_44) begin
      dl_out_data_44 <= dat_out_bypass_data_44;
    end
    if (dat_out_mask_45) begin
      dl_out_data_45 <= dat_out_bypass_data_45;
    end
    if (dat_out_mask_46) begin
      dl_out_data_46 <= dat_out_bypass_data_46;
    end
    if (dat_out_mask_47) begin
      dl_out_data_47 <= dat_out_bypass_data_47;
    end
    if (dat_out_mask_48) begin
      dl_out_data_48 <= dat_out_bypass_data_48;
    end
    if (dat_out_mask_49) begin
      dl_out_data_49 <= dat_out_bypass_data_49;
    end
    if (dat_out_mask_50) begin
      dl_out_data_50 <= dat_out_bypass_data_50;
    end
    if (dat_out_mask_51) begin
      dl_out_data_51 <= dat_out_bypass_data_51;
    end
    if (dat_out_mask_52) begin
      dl_out_data_52 <= dat_out_bypass_data_52;
    end
    if (dat_out_mask_53) begin
      dl_out_data_53 <= dat_out_bypass_data_53;
    end
    if (dat_out_mask_54) begin
      dl_out_data_54 <= dat_out_bypass_data_54;
    end
    if (dat_out_mask_55) begin
      dl_out_data_55 <= dat_out_bypass_data_55;
    end
    if (dat_out_mask_56) begin
      dl_out_data_56 <= dat_out_bypass_data_56;
    end
    if (dat_out_mask_57) begin
      dl_out_data_57 <= dat_out_bypass_data_57;
    end
    if (dat_out_mask_58) begin
      dl_out_data_58 <= dat_out_bypass_data_58;
    end
    if (dat_out_mask_59) begin
      dl_out_data_59 <= dat_out_bypass_data_59;
    end
    if (dat_out_mask_60) begin
      dl_out_data_60 <= dat_out_bypass_data_60;
    end
    if (dat_out_mask_61) begin
      dl_out_data_61 <= dat_out_bypass_data_61;
    end
    if (dat_out_mask_62) begin
      dl_out_data_62 <= dat_out_bypass_data_62;
    end
    if (dat_out_mask_63) begin
      dl_out_data_63 <= dat_out_bypass_data_63;
    end
    if (_T_337) begin
      dl_out_pvld_d1 <= 1'h0;
    end else begin
      dl_out_pvld_d1 <= dl_out_pvld;
    end
    if (_T_337) begin
      _T_4119 <= 1'h0;
    end else begin
      _T_4119 <= dl_out_pvld;
    end
    if (_T_337) begin
      _T_4122 <= 1'h0;
    end else begin
      _T_4122 <= dl_out_pvld;
    end
    if (_T_337) begin
      _T_4126 <= 9'h0;
    end else begin
      if (_T_4124) begin
        if (_T_4115) begin
          _T_4126 <= 9'h0;
        end else begin
          _T_4126 <= dl_out_flag;
        end
      end
    end
    if (_T_337) begin
      _T_4130 <= 9'h0;
    end else begin
      if (_T_4124) begin
        if (_T_4115) begin
          _T_4130 <= 9'h0;
        end else begin
          _T_4130 <= dl_out_flag;
        end
      end
    end
    if (_T_337) begin
      _T_4398_0 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_0 <= dl_out_mask_0;
      end
    end
    if (_T_337) begin
      _T_4398_1 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_1 <= dl_out_mask_1;
      end
    end
    if (_T_337) begin
      _T_4398_2 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_2 <= dl_out_mask_2;
      end
    end
    if (_T_337) begin
      _T_4398_3 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_3 <= dl_out_mask_3;
      end
    end
    if (_T_337) begin
      _T_4398_4 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_4 <= dl_out_mask_4;
      end
    end
    if (_T_337) begin
      _T_4398_5 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_5 <= dl_out_mask_5;
      end
    end
    if (_T_337) begin
      _T_4398_6 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_6 <= dl_out_mask_6;
      end
    end
    if (_T_337) begin
      _T_4398_7 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_7 <= dl_out_mask_7;
      end
    end
    if (_T_337) begin
      _T_4398_8 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_8 <= dl_out_mask_8;
      end
    end
    if (_T_337) begin
      _T_4398_9 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_9 <= dl_out_mask_9;
      end
    end
    if (_T_337) begin
      _T_4398_10 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_10 <= dl_out_mask_10;
      end
    end
    if (_T_337) begin
      _T_4398_11 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_11 <= dl_out_mask_11;
      end
    end
    if (_T_337) begin
      _T_4398_12 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_12 <= dl_out_mask_12;
      end
    end
    if (_T_337) begin
      _T_4398_13 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_13 <= dl_out_mask_13;
      end
    end
    if (_T_337) begin
      _T_4398_14 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_14 <= dl_out_mask_14;
      end
    end
    if (_T_337) begin
      _T_4398_15 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_15 <= dl_out_mask_15;
      end
    end
    if (_T_337) begin
      _T_4398_16 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_16 <= dl_out_mask_16;
      end
    end
    if (_T_337) begin
      _T_4398_17 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_17 <= dl_out_mask_17;
      end
    end
    if (_T_337) begin
      _T_4398_18 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_18 <= dl_out_mask_18;
      end
    end
    if (_T_337) begin
      _T_4398_19 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_19 <= dl_out_mask_19;
      end
    end
    if (_T_337) begin
      _T_4398_20 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_20 <= dl_out_mask_20;
      end
    end
    if (_T_337) begin
      _T_4398_21 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_21 <= dl_out_mask_21;
      end
    end
    if (_T_337) begin
      _T_4398_22 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_22 <= dl_out_mask_22;
      end
    end
    if (_T_337) begin
      _T_4398_23 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_23 <= dl_out_mask_23;
      end
    end
    if (_T_337) begin
      _T_4398_24 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_24 <= dl_out_mask_24;
      end
    end
    if (_T_337) begin
      _T_4398_25 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_25 <= dl_out_mask_25;
      end
    end
    if (_T_337) begin
      _T_4398_26 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_26 <= dl_out_mask_26;
      end
    end
    if (_T_337) begin
      _T_4398_27 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_27 <= dl_out_mask_27;
      end
    end
    if (_T_337) begin
      _T_4398_28 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_28 <= dl_out_mask_28;
      end
    end
    if (_T_337) begin
      _T_4398_29 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_29 <= dl_out_mask_29;
      end
    end
    if (_T_337) begin
      _T_4398_30 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_30 <= dl_out_mask_30;
      end
    end
    if (_T_337) begin
      _T_4398_31 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_31 <= dl_out_mask_31;
      end
    end
    if (_T_337) begin
      _T_4398_32 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_32 <= dl_out_mask_32;
      end
    end
    if (_T_337) begin
      _T_4398_33 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_33 <= dl_out_mask_33;
      end
    end
    if (_T_337) begin
      _T_4398_34 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_34 <= dl_out_mask_34;
      end
    end
    if (_T_337) begin
      _T_4398_35 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_35 <= dl_out_mask_35;
      end
    end
    if (_T_337) begin
      _T_4398_36 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_36 <= dl_out_mask_36;
      end
    end
    if (_T_337) begin
      _T_4398_37 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_37 <= dl_out_mask_37;
      end
    end
    if (_T_337) begin
      _T_4398_38 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_38 <= dl_out_mask_38;
      end
    end
    if (_T_337) begin
      _T_4398_39 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_39 <= dl_out_mask_39;
      end
    end
    if (_T_337) begin
      _T_4398_40 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_40 <= dl_out_mask_40;
      end
    end
    if (_T_337) begin
      _T_4398_41 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_41 <= dl_out_mask_41;
      end
    end
    if (_T_337) begin
      _T_4398_42 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_42 <= dl_out_mask_42;
      end
    end
    if (_T_337) begin
      _T_4398_43 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_43 <= dl_out_mask_43;
      end
    end
    if (_T_337) begin
      _T_4398_44 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_44 <= dl_out_mask_44;
      end
    end
    if (_T_337) begin
      _T_4398_45 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_45 <= dl_out_mask_45;
      end
    end
    if (_T_337) begin
      _T_4398_46 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_46 <= dl_out_mask_46;
      end
    end
    if (_T_337) begin
      _T_4398_47 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_47 <= dl_out_mask_47;
      end
    end
    if (_T_337) begin
      _T_4398_48 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_48 <= dl_out_mask_48;
      end
    end
    if (_T_337) begin
      _T_4398_49 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_49 <= dl_out_mask_49;
      end
    end
    if (_T_337) begin
      _T_4398_50 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_50 <= dl_out_mask_50;
      end
    end
    if (_T_337) begin
      _T_4398_51 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_51 <= dl_out_mask_51;
      end
    end
    if (_T_337) begin
      _T_4398_52 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_52 <= dl_out_mask_52;
      end
    end
    if (_T_337) begin
      _T_4398_53 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_53 <= dl_out_mask_53;
      end
    end
    if (_T_337) begin
      _T_4398_54 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_54 <= dl_out_mask_54;
      end
    end
    if (_T_337) begin
      _T_4398_55 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_55 <= dl_out_mask_55;
      end
    end
    if (_T_337) begin
      _T_4398_56 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_56 <= dl_out_mask_56;
      end
    end
    if (_T_337) begin
      _T_4398_57 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_57 <= dl_out_mask_57;
      end
    end
    if (_T_337) begin
      _T_4398_58 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_58 <= dl_out_mask_58;
      end
    end
    if (_T_337) begin
      _T_4398_59 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_59 <= dl_out_mask_59;
      end
    end
    if (_T_337) begin
      _T_4398_60 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_60 <= dl_out_mask_60;
      end
    end
    if (_T_337) begin
      _T_4398_61 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_61 <= dl_out_mask_61;
      end
    end
    if (_T_337) begin
      _T_4398_62 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_62 <= dl_out_mask_62;
      end
    end
    if (_T_337) begin
      _T_4398_63 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4398_63 <= dl_out_mask_63;
      end
    end
    if (_T_337) begin
      _T_4925_0 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_0 <= dl_out_mask_0;
      end
    end
    if (_T_337) begin
      _T_4925_1 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_1 <= dl_out_mask_1;
      end
    end
    if (_T_337) begin
      _T_4925_2 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_2 <= dl_out_mask_2;
      end
    end
    if (_T_337) begin
      _T_4925_3 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_3 <= dl_out_mask_3;
      end
    end
    if (_T_337) begin
      _T_4925_4 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_4 <= dl_out_mask_4;
      end
    end
    if (_T_337) begin
      _T_4925_5 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_5 <= dl_out_mask_5;
      end
    end
    if (_T_337) begin
      _T_4925_6 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_6 <= dl_out_mask_6;
      end
    end
    if (_T_337) begin
      _T_4925_7 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_7 <= dl_out_mask_7;
      end
    end
    if (_T_337) begin
      _T_4925_8 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_8 <= dl_out_mask_8;
      end
    end
    if (_T_337) begin
      _T_4925_9 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_9 <= dl_out_mask_9;
      end
    end
    if (_T_337) begin
      _T_4925_10 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_10 <= dl_out_mask_10;
      end
    end
    if (_T_337) begin
      _T_4925_11 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_11 <= dl_out_mask_11;
      end
    end
    if (_T_337) begin
      _T_4925_12 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_12 <= dl_out_mask_12;
      end
    end
    if (_T_337) begin
      _T_4925_13 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_13 <= dl_out_mask_13;
      end
    end
    if (_T_337) begin
      _T_4925_14 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_14 <= dl_out_mask_14;
      end
    end
    if (_T_337) begin
      _T_4925_15 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_15 <= dl_out_mask_15;
      end
    end
    if (_T_337) begin
      _T_4925_16 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_16 <= dl_out_mask_16;
      end
    end
    if (_T_337) begin
      _T_4925_17 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_17 <= dl_out_mask_17;
      end
    end
    if (_T_337) begin
      _T_4925_18 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_18 <= dl_out_mask_18;
      end
    end
    if (_T_337) begin
      _T_4925_19 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_19 <= dl_out_mask_19;
      end
    end
    if (_T_337) begin
      _T_4925_20 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_20 <= dl_out_mask_20;
      end
    end
    if (_T_337) begin
      _T_4925_21 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_21 <= dl_out_mask_21;
      end
    end
    if (_T_337) begin
      _T_4925_22 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_22 <= dl_out_mask_22;
      end
    end
    if (_T_337) begin
      _T_4925_23 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_23 <= dl_out_mask_23;
      end
    end
    if (_T_337) begin
      _T_4925_24 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_24 <= dl_out_mask_24;
      end
    end
    if (_T_337) begin
      _T_4925_25 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_25 <= dl_out_mask_25;
      end
    end
    if (_T_337) begin
      _T_4925_26 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_26 <= dl_out_mask_26;
      end
    end
    if (_T_337) begin
      _T_4925_27 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_27 <= dl_out_mask_27;
      end
    end
    if (_T_337) begin
      _T_4925_28 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_28 <= dl_out_mask_28;
      end
    end
    if (_T_337) begin
      _T_4925_29 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_29 <= dl_out_mask_29;
      end
    end
    if (_T_337) begin
      _T_4925_30 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_30 <= dl_out_mask_30;
      end
    end
    if (_T_337) begin
      _T_4925_31 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_31 <= dl_out_mask_31;
      end
    end
    if (_T_337) begin
      _T_4925_32 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_32 <= dl_out_mask_32;
      end
    end
    if (_T_337) begin
      _T_4925_33 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_33 <= dl_out_mask_33;
      end
    end
    if (_T_337) begin
      _T_4925_34 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_34 <= dl_out_mask_34;
      end
    end
    if (_T_337) begin
      _T_4925_35 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_35 <= dl_out_mask_35;
      end
    end
    if (_T_337) begin
      _T_4925_36 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_36 <= dl_out_mask_36;
      end
    end
    if (_T_337) begin
      _T_4925_37 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_37 <= dl_out_mask_37;
      end
    end
    if (_T_337) begin
      _T_4925_38 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_38 <= dl_out_mask_38;
      end
    end
    if (_T_337) begin
      _T_4925_39 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_39 <= dl_out_mask_39;
      end
    end
    if (_T_337) begin
      _T_4925_40 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_40 <= dl_out_mask_40;
      end
    end
    if (_T_337) begin
      _T_4925_41 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_41 <= dl_out_mask_41;
      end
    end
    if (_T_337) begin
      _T_4925_42 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_42 <= dl_out_mask_42;
      end
    end
    if (_T_337) begin
      _T_4925_43 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_43 <= dl_out_mask_43;
      end
    end
    if (_T_337) begin
      _T_4925_44 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_44 <= dl_out_mask_44;
      end
    end
    if (_T_337) begin
      _T_4925_45 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_45 <= dl_out_mask_45;
      end
    end
    if (_T_337) begin
      _T_4925_46 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_46 <= dl_out_mask_46;
      end
    end
    if (_T_337) begin
      _T_4925_47 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_47 <= dl_out_mask_47;
      end
    end
    if (_T_337) begin
      _T_4925_48 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_48 <= dl_out_mask_48;
      end
    end
    if (_T_337) begin
      _T_4925_49 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_49 <= dl_out_mask_49;
      end
    end
    if (_T_337) begin
      _T_4925_50 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_50 <= dl_out_mask_50;
      end
    end
    if (_T_337) begin
      _T_4925_51 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_51 <= dl_out_mask_51;
      end
    end
    if (_T_337) begin
      _T_4925_52 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_52 <= dl_out_mask_52;
      end
    end
    if (_T_337) begin
      _T_4925_53 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_53 <= dl_out_mask_53;
      end
    end
    if (_T_337) begin
      _T_4925_54 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_54 <= dl_out_mask_54;
      end
    end
    if (_T_337) begin
      _T_4925_55 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_55 <= dl_out_mask_55;
      end
    end
    if (_T_337) begin
      _T_4925_56 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_56 <= dl_out_mask_56;
      end
    end
    if (_T_337) begin
      _T_4925_57 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_57 <= dl_out_mask_57;
      end
    end
    if (_T_337) begin
      _T_4925_58 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_58 <= dl_out_mask_58;
      end
    end
    if (_T_337) begin
      _T_4925_59 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_59 <= dl_out_mask_59;
      end
    end
    if (_T_337) begin
      _T_4925_60 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_60 <= dl_out_mask_60;
      end
    end
    if (_T_337) begin
      _T_4925_61 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_61 <= dl_out_mask_61;
      end
    end
    if (_T_337) begin
      _T_4925_62 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_62 <= dl_out_mask_62;
      end
    end
    if (_T_337) begin
      _T_4925_63 <= 1'h0;
    end else begin
      if (_T_4124) begin
        _T_4925_63 <= dl_out_mask_63;
      end
    end
    if (dl_out_mask_0) begin
      _T_5186 <= dl_out_data_0;
    end
    if (dl_out_mask_0) begin
      _T_5188 <= dl_out_data_0;
    end
    if (dl_out_mask_1) begin
      _T_5190 <= dl_out_data_1;
    end
    if (dl_out_mask_1) begin
      _T_5192 <= dl_out_data_1;
    end
    if (dl_out_mask_2) begin
      _T_5194 <= dl_out_data_2;
    end
    if (dl_out_mask_2) begin
      _T_5196 <= dl_out_data_2;
    end
    if (dl_out_mask_3) begin
      _T_5198 <= dl_out_data_3;
    end
    if (dl_out_mask_3) begin
      _T_5200 <= dl_out_data_3;
    end
    if (dl_out_mask_4) begin
      _T_5202 <= dl_out_data_4;
    end
    if (dl_out_mask_4) begin
      _T_5204 <= dl_out_data_4;
    end
    if (dl_out_mask_5) begin
      _T_5206 <= dl_out_data_5;
    end
    if (dl_out_mask_5) begin
      _T_5208 <= dl_out_data_5;
    end
    if (dl_out_mask_6) begin
      _T_5210 <= dl_out_data_6;
    end
    if (dl_out_mask_6) begin
      _T_5212 <= dl_out_data_6;
    end
    if (dl_out_mask_7) begin
      _T_5214 <= dl_out_data_7;
    end
    if (dl_out_mask_7) begin
      _T_5216 <= dl_out_data_7;
    end
    if (dl_out_mask_8) begin
      _T_5218 <= dl_out_data_8;
    end
    if (dl_out_mask_8) begin
      _T_5220 <= dl_out_data_8;
    end
    if (dl_out_mask_9) begin
      _T_5222 <= dl_out_data_9;
    end
    if (dl_out_mask_9) begin
      _T_5224 <= dl_out_data_9;
    end
    if (dl_out_mask_10) begin
      _T_5226 <= dl_out_data_10;
    end
    if (dl_out_mask_10) begin
      _T_5228 <= dl_out_data_10;
    end
    if (dl_out_mask_11) begin
      _T_5230 <= dl_out_data_11;
    end
    if (dl_out_mask_11) begin
      _T_5232 <= dl_out_data_11;
    end
    if (dl_out_mask_12) begin
      _T_5234 <= dl_out_data_12;
    end
    if (dl_out_mask_12) begin
      _T_5236 <= dl_out_data_12;
    end
    if (dl_out_mask_13) begin
      _T_5238 <= dl_out_data_13;
    end
    if (dl_out_mask_13) begin
      _T_5240 <= dl_out_data_13;
    end
    if (dl_out_mask_14) begin
      _T_5242 <= dl_out_data_14;
    end
    if (dl_out_mask_14) begin
      _T_5244 <= dl_out_data_14;
    end
    if (dl_out_mask_15) begin
      _T_5246 <= dl_out_data_15;
    end
    if (dl_out_mask_15) begin
      _T_5248 <= dl_out_data_15;
    end
    if (dl_out_mask_16) begin
      _T_5250 <= dl_out_data_16;
    end
    if (dl_out_mask_16) begin
      _T_5252 <= dl_out_data_16;
    end
    if (dl_out_mask_17) begin
      _T_5254 <= dl_out_data_17;
    end
    if (dl_out_mask_17) begin
      _T_5256 <= dl_out_data_17;
    end
    if (dl_out_mask_18) begin
      _T_5258 <= dl_out_data_18;
    end
    if (dl_out_mask_18) begin
      _T_5260 <= dl_out_data_18;
    end
    if (dl_out_mask_19) begin
      _T_5262 <= dl_out_data_19;
    end
    if (dl_out_mask_19) begin
      _T_5264 <= dl_out_data_19;
    end
    if (dl_out_mask_20) begin
      _T_5266 <= dl_out_data_20;
    end
    if (dl_out_mask_20) begin
      _T_5268 <= dl_out_data_20;
    end
    if (dl_out_mask_21) begin
      _T_5270 <= dl_out_data_21;
    end
    if (dl_out_mask_21) begin
      _T_5272 <= dl_out_data_21;
    end
    if (dl_out_mask_22) begin
      _T_5274 <= dl_out_data_22;
    end
    if (dl_out_mask_22) begin
      _T_5276 <= dl_out_data_22;
    end
    if (dl_out_mask_23) begin
      _T_5278 <= dl_out_data_23;
    end
    if (dl_out_mask_23) begin
      _T_5280 <= dl_out_data_23;
    end
    if (dl_out_mask_24) begin
      _T_5282 <= dl_out_data_24;
    end
    if (dl_out_mask_24) begin
      _T_5284 <= dl_out_data_24;
    end
    if (dl_out_mask_25) begin
      _T_5286 <= dl_out_data_25;
    end
    if (dl_out_mask_25) begin
      _T_5288 <= dl_out_data_25;
    end
    if (dl_out_mask_26) begin
      _T_5290 <= dl_out_data_26;
    end
    if (dl_out_mask_26) begin
      _T_5292 <= dl_out_data_26;
    end
    if (dl_out_mask_27) begin
      _T_5294 <= dl_out_data_27;
    end
    if (dl_out_mask_27) begin
      _T_5296 <= dl_out_data_27;
    end
    if (dl_out_mask_28) begin
      _T_5298 <= dl_out_data_28;
    end
    if (dl_out_mask_28) begin
      _T_5300 <= dl_out_data_28;
    end
    if (dl_out_mask_29) begin
      _T_5302 <= dl_out_data_29;
    end
    if (dl_out_mask_29) begin
      _T_5304 <= dl_out_data_29;
    end
    if (dl_out_mask_30) begin
      _T_5306 <= dl_out_data_30;
    end
    if (dl_out_mask_30) begin
      _T_5308 <= dl_out_data_30;
    end
    if (dl_out_mask_31) begin
      _T_5310 <= dl_out_data_31;
    end
    if (dl_out_mask_31) begin
      _T_5312 <= dl_out_data_31;
    end
    if (dl_out_mask_32) begin
      _T_5314 <= dl_out_data_32;
    end
    if (dl_out_mask_32) begin
      _T_5316 <= dl_out_data_32;
    end
    if (dl_out_mask_33) begin
      _T_5318 <= dl_out_data_33;
    end
    if (dl_out_mask_33) begin
      _T_5320 <= dl_out_data_33;
    end
    if (dl_out_mask_34) begin
      _T_5322 <= dl_out_data_34;
    end
    if (dl_out_mask_34) begin
      _T_5324 <= dl_out_data_34;
    end
    if (dl_out_mask_35) begin
      _T_5326 <= dl_out_data_35;
    end
    if (dl_out_mask_35) begin
      _T_5328 <= dl_out_data_35;
    end
    if (dl_out_mask_36) begin
      _T_5330 <= dl_out_data_36;
    end
    if (dl_out_mask_36) begin
      _T_5332 <= dl_out_data_36;
    end
    if (dl_out_mask_37) begin
      _T_5334 <= dl_out_data_37;
    end
    if (dl_out_mask_37) begin
      _T_5336 <= dl_out_data_37;
    end
    if (dl_out_mask_38) begin
      _T_5338 <= dl_out_data_38;
    end
    if (dl_out_mask_38) begin
      _T_5340 <= dl_out_data_38;
    end
    if (dl_out_mask_39) begin
      _T_5342 <= dl_out_data_39;
    end
    if (dl_out_mask_39) begin
      _T_5344 <= dl_out_data_39;
    end
    if (dl_out_mask_40) begin
      _T_5346 <= dl_out_data_40;
    end
    if (dl_out_mask_40) begin
      _T_5348 <= dl_out_data_40;
    end
    if (dl_out_mask_41) begin
      _T_5350 <= dl_out_data_41;
    end
    if (dl_out_mask_41) begin
      _T_5352 <= dl_out_data_41;
    end
    if (dl_out_mask_42) begin
      _T_5354 <= dl_out_data_42;
    end
    if (dl_out_mask_42) begin
      _T_5356 <= dl_out_data_42;
    end
    if (dl_out_mask_43) begin
      _T_5358 <= dl_out_data_43;
    end
    if (dl_out_mask_43) begin
      _T_5360 <= dl_out_data_43;
    end
    if (dl_out_mask_44) begin
      _T_5362 <= dl_out_data_44;
    end
    if (dl_out_mask_44) begin
      _T_5364 <= dl_out_data_44;
    end
    if (dl_out_mask_45) begin
      _T_5366 <= dl_out_data_45;
    end
    if (dl_out_mask_45) begin
      _T_5368 <= dl_out_data_45;
    end
    if (dl_out_mask_46) begin
      _T_5370 <= dl_out_data_46;
    end
    if (dl_out_mask_46) begin
      _T_5372 <= dl_out_data_46;
    end
    if (dl_out_mask_47) begin
      _T_5374 <= dl_out_data_47;
    end
    if (dl_out_mask_47) begin
      _T_5376 <= dl_out_data_47;
    end
    if (dl_out_mask_48) begin
      _T_5378 <= dl_out_data_48;
    end
    if (dl_out_mask_48) begin
      _T_5380 <= dl_out_data_48;
    end
    if (dl_out_mask_49) begin
      _T_5382 <= dl_out_data_49;
    end
    if (dl_out_mask_49) begin
      _T_5384 <= dl_out_data_49;
    end
    if (dl_out_mask_50) begin
      _T_5386 <= dl_out_data_50;
    end
    if (dl_out_mask_50) begin
      _T_5388 <= dl_out_data_50;
    end
    if (dl_out_mask_51) begin
      _T_5390 <= dl_out_data_51;
    end
    if (dl_out_mask_51) begin
      _T_5392 <= dl_out_data_51;
    end
    if (dl_out_mask_52) begin
      _T_5394 <= dl_out_data_52;
    end
    if (dl_out_mask_52) begin
      _T_5396 <= dl_out_data_52;
    end
    if (dl_out_mask_53) begin
      _T_5398 <= dl_out_data_53;
    end
    if (dl_out_mask_53) begin
      _T_5400 <= dl_out_data_53;
    end
    if (dl_out_mask_54) begin
      _T_5402 <= dl_out_data_54;
    end
    if (dl_out_mask_54) begin
      _T_5404 <= dl_out_data_54;
    end
    if (dl_out_mask_55) begin
      _T_5406 <= dl_out_data_55;
    end
    if (dl_out_mask_55) begin
      _T_5408 <= dl_out_data_55;
    end
    if (dl_out_mask_56) begin
      _T_5410 <= dl_out_data_56;
    end
    if (dl_out_mask_56) begin
      _T_5412 <= dl_out_data_56;
    end
    if (dl_out_mask_57) begin
      _T_5414 <= dl_out_data_57;
    end
    if (dl_out_mask_57) begin
      _T_5416 <= dl_out_data_57;
    end
    if (dl_out_mask_58) begin
      _T_5418 <= dl_out_data_58;
    end
    if (dl_out_mask_58) begin
      _T_5420 <= dl_out_data_58;
    end
    if (dl_out_mask_59) begin
      _T_5422 <= dl_out_data_59;
    end
    if (dl_out_mask_59) begin
      _T_5424 <= dl_out_data_59;
    end
    if (dl_out_mask_60) begin
      _T_5426 <= dl_out_data_60;
    end
    if (dl_out_mask_60) begin
      _T_5428 <= dl_out_data_60;
    end
    if (dl_out_mask_61) begin
      _T_5430 <= dl_out_data_61;
    end
    if (dl_out_mask_61) begin
      _T_5432 <= dl_out_data_61;
    end
    if (dl_out_mask_62) begin
      _T_5434 <= dl_out_data_62;
    end
    if (dl_out_mask_62) begin
      _T_5436 <= dl_out_data_62;
    end
    if (dl_out_mask_63) begin
      _T_5438 <= dl_out_data_63;
    end
    if (dl_out_mask_63) begin
      _T_5440 <= dl_out_data_63;
    end
  end
  always @(posedge nvdla_core_ng_clk) begin
    if (_T_337) begin
      dat_entry_st <= 15'h0;
    end else begin
      if (_T_758) begin
        if (sc2cdma_dat_pending_req) begin
          dat_entry_st <= 15'h0;
        end else begin
          if (is_dat_entry_st_wrap) begin
            dat_entry_st <= dat_entry_st_inc_wrap;
          end else begin
            dat_entry_st <= dat_entry_st_inc;
          end
        end
      end
    end
  end
endmodule



// ================================================================
// NVDLA Open Source Project
//
// Copyright(c) 2016 - 2017 NVIDIA Corporation. Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CSC_dl.v
// ================================================================
// NVDLA Open Source Project
// 
// Copyright(c) 2016 - 2017 NVIDIA Corporation.  Licensed under the
// NVDLA Open Hardware License; Check "LICENSE" which comes with 
// this distribution for more information.
// ================================================================
// File Name: NV_NVDLA_CSC.h

module NV_NVDLA_CSC_dl (
   nvdla_core_clk //|< i
  ,nvdla_core_rstn //|< i
  ,sg2dl_pvld //|< i
  ,sg2dl_pd //|< i
  ,sc_state //|< i
  ,sg2dl_reuse_rls //|< i
  ,sc2cdma_dat_pending_req //|< i
  ,cdma2sc_dat_updt //|< i
  ,cdma2sc_dat_entries //|< i
  ,cdma2sc_dat_slices //|< i
  ,sc2cdma_dat_updt //|> o
  ,sc2cdma_dat_entries //|> o
  ,sc2cdma_dat_slices //|> o
  ,sc2buf_dat_rd_en //|> o
  ,sc2buf_dat_rd_addr //|> o
  ,sc2buf_dat_rd_valid //|< i
  ,sc2buf_dat_rd_data //|< i
  ,sc2mac_dat_a_pvld //|> o
  ,sc2mac_dat_a_mask //|> o
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: ,sc2mac_dat_a_data${i} //|> o )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,sc2mac_dat_a_data0 //|> o 
,sc2mac_dat_a_data1 //|> o 
,sc2mac_dat_a_data2 //|> o 
,sc2mac_dat_a_data3 //|> o 
,sc2mac_dat_a_data4 //|> o 
,sc2mac_dat_a_data5 //|> o 
,sc2mac_dat_a_data6 //|> o 
,sc2mac_dat_a_data7 //|> o 
,sc2mac_dat_a_data8 //|> o 
,sc2mac_dat_a_data9 //|> o 
,sc2mac_dat_a_data10 //|> o 
,sc2mac_dat_a_data11 //|> o 
,sc2mac_dat_a_data12 //|> o 
,sc2mac_dat_a_data13 //|> o 
,sc2mac_dat_a_data14 //|> o 
,sc2mac_dat_a_data15 //|> o 
,sc2mac_dat_a_data16 //|> o 
,sc2mac_dat_a_data17 //|> o 
,sc2mac_dat_a_data18 //|> o 
,sc2mac_dat_a_data19 //|> o 
,sc2mac_dat_a_data20 //|> o 
,sc2mac_dat_a_data21 //|> o 
,sc2mac_dat_a_data22 //|> o 
,sc2mac_dat_a_data23 //|> o 
,sc2mac_dat_a_data24 //|> o 
,sc2mac_dat_a_data25 //|> o 
,sc2mac_dat_a_data26 //|> o 
,sc2mac_dat_a_data27 //|> o 
,sc2mac_dat_a_data28 //|> o 
,sc2mac_dat_a_data29 //|> o 
,sc2mac_dat_a_data30 //|> o 
,sc2mac_dat_a_data31 //|> o 
,sc2mac_dat_a_data32 //|> o 
,sc2mac_dat_a_data33 //|> o 
,sc2mac_dat_a_data34 //|> o 
,sc2mac_dat_a_data35 //|> o 
,sc2mac_dat_a_data36 //|> o 
,sc2mac_dat_a_data37 //|> o 
,sc2mac_dat_a_data38 //|> o 
,sc2mac_dat_a_data39 //|> o 
,sc2mac_dat_a_data40 //|> o 
,sc2mac_dat_a_data41 //|> o 
,sc2mac_dat_a_data42 //|> o 
,sc2mac_dat_a_data43 //|> o 
,sc2mac_dat_a_data44 //|> o 
,sc2mac_dat_a_data45 //|> o 
,sc2mac_dat_a_data46 //|> o 
,sc2mac_dat_a_data47 //|> o 
,sc2mac_dat_a_data48 //|> o 
,sc2mac_dat_a_data49 //|> o 
,sc2mac_dat_a_data50 //|> o 
,sc2mac_dat_a_data51 //|> o 
,sc2mac_dat_a_data52 //|> o 
,sc2mac_dat_a_data53 //|> o 
,sc2mac_dat_a_data54 //|> o 
,sc2mac_dat_a_data55 //|> o 
,sc2mac_dat_a_data56 //|> o 
,sc2mac_dat_a_data57 //|> o 
,sc2mac_dat_a_data58 //|> o 
,sc2mac_dat_a_data59 //|> o 
,sc2mac_dat_a_data60 //|> o 
,sc2mac_dat_a_data61 //|> o 
,sc2mac_dat_a_data62 //|> o 
,sc2mac_dat_a_data63 //|> o 
//| eperl: generated_end (DO NOT EDIT ABOVE)
  ,sc2mac_dat_a_pd //|> o
  ,sc2mac_dat_b_pvld //|> o
  ,sc2mac_dat_b_mask //|> o
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: ,sc2mac_dat_b_data${i} //|> o )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

,sc2mac_dat_b_data0 //|> o 
,sc2mac_dat_b_data1 //|> o 
,sc2mac_dat_b_data2 //|> o 
,sc2mac_dat_b_data3 //|> o 
,sc2mac_dat_b_data4 //|> o 
,sc2mac_dat_b_data5 //|> o 
,sc2mac_dat_b_data6 //|> o 
,sc2mac_dat_b_data7 //|> o 
,sc2mac_dat_b_data8 //|> o 
,sc2mac_dat_b_data9 //|> o 
,sc2mac_dat_b_data10 //|> o 
,sc2mac_dat_b_data11 //|> o 
,sc2mac_dat_b_data12 //|> o 
,sc2mac_dat_b_data13 //|> o 
,sc2mac_dat_b_data14 //|> o 
,sc2mac_dat_b_data15 //|> o 
,sc2mac_dat_b_data16 //|> o 
,sc2mac_dat_b_data17 //|> o 
,sc2mac_dat_b_data18 //|> o 
,sc2mac_dat_b_data19 //|> o 
,sc2mac_dat_b_data20 //|> o 
,sc2mac_dat_b_data21 //|> o 
,sc2mac_dat_b_data22 //|> o 
,sc2mac_dat_b_data23 //|> o 
,sc2mac_dat_b_data24 //|> o 
,sc2mac_dat_b_data25 //|> o 
,sc2mac_dat_b_data26 //|> o 
,sc2mac_dat_b_data27 //|> o 
,sc2mac_dat_b_data28 //|> o 
,sc2mac_dat_b_data29 //|> o 
,sc2mac_dat_b_data30 //|> o 
,sc2mac_dat_b_data31 //|> o 
,sc2mac_dat_b_data32 //|> o 
,sc2mac_dat_b_data33 //|> o 
,sc2mac_dat_b_data34 //|> o 
,sc2mac_dat_b_data35 //|> o 
,sc2mac_dat_b_data36 //|> o 
,sc2mac_dat_b_data37 //|> o 
,sc2mac_dat_b_data38 //|> o 
,sc2mac_dat_b_data39 //|> o 
,sc2mac_dat_b_data40 //|> o 
,sc2mac_dat_b_data41 //|> o 
,sc2mac_dat_b_data42 //|> o 
,sc2mac_dat_b_data43 //|> o 
,sc2mac_dat_b_data44 //|> o 
,sc2mac_dat_b_data45 //|> o 
,sc2mac_dat_b_data46 //|> o 
,sc2mac_dat_b_data47 //|> o 
,sc2mac_dat_b_data48 //|> o 
,sc2mac_dat_b_data49 //|> o 
,sc2mac_dat_b_data50 //|> o 
,sc2mac_dat_b_data51 //|> o 
,sc2mac_dat_b_data52 //|> o 
,sc2mac_dat_b_data53 //|> o 
,sc2mac_dat_b_data54 //|> o 
,sc2mac_dat_b_data55 //|> o 
,sc2mac_dat_b_data56 //|> o 
,sc2mac_dat_b_data57 //|> o 
,sc2mac_dat_b_data58 //|> o 
,sc2mac_dat_b_data59 //|> o 
,sc2mac_dat_b_data60 //|> o 
,sc2mac_dat_b_data61 //|> o 
,sc2mac_dat_b_data62 //|> o 
,sc2mac_dat_b_data63 //|> o 
//| eperl: generated_end (DO NOT EDIT ABOVE)
  ,sc2mac_dat_b_pd //|> o
  ,nvdla_core_ng_clk //|< i
  ,reg2dp_op_en //|< i
  ,reg2dp_conv_mode //|< i
  ,reg2dp_batches //|< i
  ,reg2dp_proc_precision //|< i
  ,reg2dp_datain_format //|< i
  ,reg2dp_skip_data_rls //|< i
  ,reg2dp_datain_channel_ext //|< i
  ,reg2dp_datain_height_ext //|< i
  ,reg2dp_datain_width_ext //|< i
  ,reg2dp_y_extension //|< i
  ,reg2dp_weight_channel_ext //|< i
  ,reg2dp_entries //|< i
  ,reg2dp_dataout_width //|< i
  ,reg2dp_rls_slices //|< i
  ,reg2dp_conv_x_stride_ext //|< i
  ,reg2dp_conv_y_stride_ext //|< i
  ,reg2dp_x_dilation_ext //|< i
  ,reg2dp_y_dilation_ext //|< i
  ,reg2dp_pad_left //|< i
  ,reg2dp_pad_top //|< i
  ,reg2dp_pad_value //|< i
  ,reg2dp_data_bank //|< i
  ,reg2dp_pra_truncate //|< i
  ,slcg_wg_en //|> o
  );
input nvdla_core_clk;
input nvdla_core_rstn;
input sg2dl_pvld; /* data valid */
input [30:0] sg2dl_pd;
input [1:0] sc_state;
input sg2dl_reuse_rls;
input sc2cdma_dat_pending_req;
input cdma2sc_dat_updt; /* data valid */
input [15 -1:0] cdma2sc_dat_entries;
input [13:0] cdma2sc_dat_slices;
output sc2cdma_dat_updt; /* data valid */
output [15 -1:0] sc2cdma_dat_entries;
output [13:0] sc2cdma_dat_slices;
output sc2buf_dat_rd_en; /* data valid */
output [13 -1:0] sc2buf_dat_rd_addr;
input sc2buf_dat_rd_valid; /* data valid */
input [512 -1:0] sc2buf_dat_rd_data;
output sc2mac_dat_a_pvld; /* data valid */
output [64 -1:0] sc2mac_dat_a_mask;
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: output [8 -1:0] sc2mac_dat_a_data${i}; )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

output [8 -1:0] sc2mac_dat_a_data0; 
output [8 -1:0] sc2mac_dat_a_data1; 
output [8 -1:0] sc2mac_dat_a_data2; 
output [8 -1:0] sc2mac_dat_a_data3; 
output [8 -1:0] sc2mac_dat_a_data4; 
output [8 -1:0] sc2mac_dat_a_data5; 
output [8 -1:0] sc2mac_dat_a_data6; 
output [8 -1:0] sc2mac_dat_a_data7; 
output [8 -1:0] sc2mac_dat_a_data8; 
output [8 -1:0] sc2mac_dat_a_data9; 
output [8 -1:0] sc2mac_dat_a_data10; 
output [8 -1:0] sc2mac_dat_a_data11; 
output [8 -1:0] sc2mac_dat_a_data12; 
output [8 -1:0] sc2mac_dat_a_data13; 
output [8 -1:0] sc2mac_dat_a_data14; 
output [8 -1:0] sc2mac_dat_a_data15; 
output [8 -1:0] sc2mac_dat_a_data16; 
output [8 -1:0] sc2mac_dat_a_data17; 
output [8 -1:0] sc2mac_dat_a_data18; 
output [8 -1:0] sc2mac_dat_a_data19; 
output [8 -1:0] sc2mac_dat_a_data20; 
output [8 -1:0] sc2mac_dat_a_data21; 
output [8 -1:0] sc2mac_dat_a_data22; 
output [8 -1:0] sc2mac_dat_a_data23; 
output [8 -1:0] sc2mac_dat_a_data24; 
output [8 -1:0] sc2mac_dat_a_data25; 
output [8 -1:0] sc2mac_dat_a_data26; 
output [8 -1:0] sc2mac_dat_a_data27; 
output [8 -1:0] sc2mac_dat_a_data28; 
output [8 -1:0] sc2mac_dat_a_data29; 
output [8 -1:0] sc2mac_dat_a_data30; 
output [8 -1:0] sc2mac_dat_a_data31; 
output [8 -1:0] sc2mac_dat_a_data32; 
output [8 -1:0] sc2mac_dat_a_data33; 
output [8 -1:0] sc2mac_dat_a_data34; 
output [8 -1:0] sc2mac_dat_a_data35; 
output [8 -1:0] sc2mac_dat_a_data36; 
output [8 -1:0] sc2mac_dat_a_data37; 
output [8 -1:0] sc2mac_dat_a_data38; 
output [8 -1:0] sc2mac_dat_a_data39; 
output [8 -1:0] sc2mac_dat_a_data40; 
output [8 -1:0] sc2mac_dat_a_data41; 
output [8 -1:0] sc2mac_dat_a_data42; 
output [8 -1:0] sc2mac_dat_a_data43; 
output [8 -1:0] sc2mac_dat_a_data44; 
output [8 -1:0] sc2mac_dat_a_data45; 
output [8 -1:0] sc2mac_dat_a_data46; 
output [8 -1:0] sc2mac_dat_a_data47; 
output [8 -1:0] sc2mac_dat_a_data48; 
output [8 -1:0] sc2mac_dat_a_data49; 
output [8 -1:0] sc2mac_dat_a_data50; 
output [8 -1:0] sc2mac_dat_a_data51; 
output [8 -1:0] sc2mac_dat_a_data52; 
output [8 -1:0] sc2mac_dat_a_data53; 
output [8 -1:0] sc2mac_dat_a_data54; 
output [8 -1:0] sc2mac_dat_a_data55; 
output [8 -1:0] sc2mac_dat_a_data56; 
output [8 -1:0] sc2mac_dat_a_data57; 
output [8 -1:0] sc2mac_dat_a_data58; 
output [8 -1:0] sc2mac_dat_a_data59; 
output [8 -1:0] sc2mac_dat_a_data60; 
output [8 -1:0] sc2mac_dat_a_data61; 
output [8 -1:0] sc2mac_dat_a_data62; 
output [8 -1:0] sc2mac_dat_a_data63; 
//| eperl: generated_end (DO NOT EDIT ABOVE)
output [8:0] sc2mac_dat_a_pd;
output sc2mac_dat_b_pvld; /* data valid */
output [64 -1:0] sc2mac_dat_b_mask;
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: output [8 -1:0] sc2mac_dat_b_data${i}; )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

output [8 -1:0] sc2mac_dat_b_data0; 
output [8 -1:0] sc2mac_dat_b_data1; 
output [8 -1:0] sc2mac_dat_b_data2; 
output [8 -1:0] sc2mac_dat_b_data3; 
output [8 -1:0] sc2mac_dat_b_data4; 
output [8 -1:0] sc2mac_dat_b_data5; 
output [8 -1:0] sc2mac_dat_b_data6; 
output [8 -1:0] sc2mac_dat_b_data7; 
output [8 -1:0] sc2mac_dat_b_data8; 
output [8 -1:0] sc2mac_dat_b_data9; 
output [8 -1:0] sc2mac_dat_b_data10; 
output [8 -1:0] sc2mac_dat_b_data11; 
output [8 -1:0] sc2mac_dat_b_data12; 
output [8 -1:0] sc2mac_dat_b_data13; 
output [8 -1:0] sc2mac_dat_b_data14; 
output [8 -1:0] sc2mac_dat_b_data15; 
output [8 -1:0] sc2mac_dat_b_data16; 
output [8 -1:0] sc2mac_dat_b_data17; 
output [8 -1:0] sc2mac_dat_b_data18; 
output [8 -1:0] sc2mac_dat_b_data19; 
output [8 -1:0] sc2mac_dat_b_data20; 
output [8 -1:0] sc2mac_dat_b_data21; 
output [8 -1:0] sc2mac_dat_b_data22; 
output [8 -1:0] sc2mac_dat_b_data23; 
output [8 -1:0] sc2mac_dat_b_data24; 
output [8 -1:0] sc2mac_dat_b_data25; 
output [8 -1:0] sc2mac_dat_b_data26; 
output [8 -1:0] sc2mac_dat_b_data27; 
output [8 -1:0] sc2mac_dat_b_data28; 
output [8 -1:0] sc2mac_dat_b_data29; 
output [8 -1:0] sc2mac_dat_b_data30; 
output [8 -1:0] sc2mac_dat_b_data31; 
output [8 -1:0] sc2mac_dat_b_data32; 
output [8 -1:0] sc2mac_dat_b_data33; 
output [8 -1:0] sc2mac_dat_b_data34; 
output [8 -1:0] sc2mac_dat_b_data35; 
output [8 -1:0] sc2mac_dat_b_data36; 
output [8 -1:0] sc2mac_dat_b_data37; 
output [8 -1:0] sc2mac_dat_b_data38; 
output [8 -1:0] sc2mac_dat_b_data39; 
output [8 -1:0] sc2mac_dat_b_data40; 
output [8 -1:0] sc2mac_dat_b_data41; 
output [8 -1:0] sc2mac_dat_b_data42; 
output [8 -1:0] sc2mac_dat_b_data43; 
output [8 -1:0] sc2mac_dat_b_data44; 
output [8 -1:0] sc2mac_dat_b_data45; 
output [8 -1:0] sc2mac_dat_b_data46; 
output [8 -1:0] sc2mac_dat_b_data47; 
output [8 -1:0] sc2mac_dat_b_data48; 
output [8 -1:0] sc2mac_dat_b_data49; 
output [8 -1:0] sc2mac_dat_b_data50; 
output [8 -1:0] sc2mac_dat_b_data51; 
output [8 -1:0] sc2mac_dat_b_data52; 
output [8 -1:0] sc2mac_dat_b_data53; 
output [8 -1:0] sc2mac_dat_b_data54; 
output [8 -1:0] sc2mac_dat_b_data55; 
output [8 -1:0] sc2mac_dat_b_data56; 
output [8 -1:0] sc2mac_dat_b_data57; 
output [8 -1:0] sc2mac_dat_b_data58; 
output [8 -1:0] sc2mac_dat_b_data59; 
output [8 -1:0] sc2mac_dat_b_data60; 
output [8 -1:0] sc2mac_dat_b_data61; 
output [8 -1:0] sc2mac_dat_b_data62; 
output [8 -1:0] sc2mac_dat_b_data63; 
//| eperl: generated_end (DO NOT EDIT ABOVE)
output [8:0] sc2mac_dat_b_pd;
input nvdla_core_ng_clk;
input [0:0] reg2dp_op_en;
input [0:0] reg2dp_conv_mode;
input [4:0] reg2dp_batches;
input [1:0] reg2dp_proc_precision;
input [0:0] reg2dp_datain_format;
input [0:0] reg2dp_skip_data_rls;
input [12:0] reg2dp_datain_channel_ext;
input [12:0] reg2dp_datain_height_ext;
input [12:0] reg2dp_datain_width_ext;
input [1:0] reg2dp_y_extension;
input [12:0] reg2dp_weight_channel_ext;
input [13:0] reg2dp_entries;
input [12:0] reg2dp_dataout_width;
input [11:0] reg2dp_rls_slices;
input [2:0] reg2dp_conv_x_stride_ext;
input [2:0] reg2dp_conv_y_stride_ext;
input [4:0] reg2dp_x_dilation_ext;
input [4:0] reg2dp_y_dilation_ext;
input [4:0] reg2dp_pad_left;
input [4:0] reg2dp_pad_top;
input [15:0] reg2dp_pad_value;
input [4:0] reg2dp_data_bank;
input [1:0] reg2dp_pra_truncate;
output slcg_wg_en;
reg [4:0] batch_cmp;
reg [4:0] batch_cnt;
reg [13 -1:0] c_bias;
reg [13 -1:0] c_bias_d1;
reg [3:0] conv_x_stride;
reg [3:0] conv_y_stride;
reg [15 -1:0] dat_entry_avl;
reg [15 -1:0] dat_entry_end;
reg [15 -1:0] dat_entry_st;
reg dat_exec_valid_d1;
reg dat_exec_valid_d2;
reg dat_l0c0_dummy;
reg [512 -1:0] dat_l0c0;
reg dat_l0c1_dummy;
reg [512 -1:0] dat_l0c1;
reg dat_l1c0_dummy;
reg [512 -1:0] dat_l1c0;
reg dat_l1c1_dummy;
reg [512 -1:0] dat_l1c1;
reg dat_l2c0_dummy;
reg [512 -1:0] dat_l2c0;
reg dat_l2c1_dummy;
reg [512 -1:0] dat_l2c1;
reg dat_l3c0_dummy;
reg [512 -1:0] dat_l3c0;
reg dat_l3c1_dummy;
reg [512 -1:0] dat_l3c1;
reg [512 -1:0] dat_out_bypass_data;
reg [64 -1:0] dat_out_bypass_mask;
reg [8:0] dat_out_flag;
reg dat_out_pvld;
reg dat_pipe_local_valid;
reg dat_pipe_valid_d1;
reg dat_pipe_valid_d2;
reg [7:0] dat_req_bytes_d1;
reg [7:0] dat_req_bytes_d2;
reg dat_req_ch_end_d1;
reg dat_req_ch_end_d2;
reg [1:0] dat_req_cur_sub_h_d1;
reg [1:0] dat_req_cur_sub_h_d2;
reg dat_req_dummy_d1;
reg dat_req_dummy_d2;
reg [8:0] dat_req_flag_d1;
reg [8:0] dat_req_flag_d2;
reg dat_req_rls_d1;
reg dat_req_rls_d2;
reg dat_req_sub_c_d1;
reg dat_req_sub_c_d2;
reg [13 -1:0] dat_req_sub_h_0_addr;
reg [13 -1:0] dat_req_sub_h_1_addr;
reg [13 -1:0] dat_req_sub_h_2_addr;
reg [13 -1:0] dat_req_sub_h_3_addr;
reg [1:0] dat_req_sub_h_d1;
reg [1:0] dat_req_sub_h_d2;
reg [1:0] dat_req_sub_w_d1;
reg [1:0] dat_req_sub_w_d2;
reg dat_req_sub_w_st_d1;
reg dat_req_sub_w_st_d2;
reg dat_req_valid_d1;
wire [512 -1:0] dat_rsp_l0_sft;
reg [512 -1:0] dat_rsp_l0_sft_d1;
reg [512 -1:0] dat_rsp_l0_sft_d2;
reg [512 -1:0] dat_rsp_l0_sft_d3;
wire [512 -1:0] dat_rsp_l1_sft;
reg [512 -1:0] dat_rsp_l1_sft_d2;
reg [512 -1:0] dat_rsp_l1_sft_d3;
wire [512 -1:0] dat_rsp_l2_sft;
reg [512 -1:0] dat_rsp_l2_sft_d3;
wire [512 -1:0] dat_rsp_l3_sft;
reg [26:0] dat_rsp_pd_d1;
reg [26:0] dat_rsp_pd_d2;
reg [26:0] dat_rsp_pd_d3;
reg [26:0] dat_rsp_pd_d4;
reg [3:0] dat_rsp_pra_en_d1;
reg dat_rsp_pvld_d1;
reg dat_rsp_pvld_d2;
reg dat_rsp_pvld_d3;
reg dat_rsp_pvld_d4;
reg [255:0] dat_rsp_wg_ch0_d1;
reg [255:0] dat_rsp_wg_ch1_d1;
reg [255:0] dat_rsp_wg_ch2_d1;
reg [255:0] dat_rsp_wg_ch3_d1;
reg [13:0] dat_slice_avl;
reg [4:0] data_bank;
reg [5:0] data_batch;
reg [10:0] datain_c_cnt;
reg [10:0] datain_channel_cmp;
reg [13:0] datain_h_cnt;
reg [13:0] datain_h_ori;
reg [12:0] datain_height_cmp;
reg [13:0] datain_w_cnt;
reg [13:0] datain_w_ori;
reg [13:0] datain_width;
reg [12:0] datain_width_cmp;
reg [12:0] dataout_w_cnt;
reg [12:0] dataout_w_ori;
reg [12:0] dataout_width_cmp;
reg [8:0] dl_out_flag;
reg [64 -1:0] dl_out_mask;
reg dl_out_pvld;
reg dl_out_pvld_d1;
reg [30:0] dl_pd_d1;
reg [30:0] dl_pd_d2;
reg [30:0] dl_pd_d3;
reg [30:0] dl_pd_d4;
reg dl_pvld_d1;
reg dl_pvld_d2;
reg dl_pvld_d3;
reg dl_pvld_d4;
reg [15 -1:0] entries;
reg [15 -1:0] entries_batch;
reg [15 -1:0] entries_cmp;
reg [13 -1:0] h_bias_0_d1;
reg [13 -1:0] h_bias_0_stride;
reg [13 -1:0] h_bias_1_d1;
reg [13 -1:0] h_bias_1_stride;
reg [13 -1:0] h_bias_2_d1;
reg [13 -1:0] h_bias_2_stride;
reg [13 -1:0] h_bias_3_d1;
reg [13 -1:0] h_bias_3_stride;
reg [13:0] h_offset_slice;
reg [33:0] is_img_d1;
reg is_sg_running_d1;
reg [21:0] is_winograd_d1;
reg [15 -1:0] last_entries;
reg [13:0] last_slices;
reg layer_st_d1;
reg [15:0] pad_value;
reg [11:0] pixel_ch_stride;
reg pixel_force_clr_d1;
reg pixel_force_fetch_d1;
reg [15:0] pixel_w_ch_ori;
reg [15:0] pixel_w_cnt;
reg [15:0] pixel_w_ori;
reg [6:0] pixel_x_add;
reg [6:0] pixel_x_byte_stride;
reg [5:0] pixel_x_init;
reg [6:0] pixel_x_init_offset;
reg pixel_x_stride_odd;
reg [7:0] pra_precision;
reg [7:0] pra_truncate;
reg [15 -1:0] rls_entries;
reg [13:0] rls_slices;
reg [7:0] rsp_sft_cnt_l0;
reg [7:0] rsp_sft_cnt_l0_ori;
reg [7:0] rsp_sft_cnt_l1;
reg [7:0] rsp_sft_cnt_l1_ori;
reg [7:0] rsp_sft_cnt_l2;
reg [7:0] rsp_sft_cnt_l2_ori;
reg [7:0] rsp_sft_cnt_l3;
reg [7:0] rsp_sft_cnt_l3_ori;
reg [13 -1:0] sc2buf_dat_rd_addr;
reg [13 -1:0] sc2buf_dat_rd_next1_addr;
reg sc2buf_dat_rd_en;
reg [15 -1:0] sc2cdma_dat_entries;
reg [13:0] sc2cdma_dat_slices;
reg sc2cdma_dat_updt;
reg [64 -1:0] sc2mac_dat_a_mask;
reg [8:0] sc2mac_dat_a_pd;
reg sc2mac_dat_a_pvld;
reg [64 -1:0] sc2mac_dat_b_mask;
reg [8:0] sc2mac_dat_b_pd;
reg sc2mac_dat_b_pvld;
reg slcg_wg_en_d1;
reg slcg_wg_en_d2;
reg slcg_wg_en_d3;
reg [13:0] slice_left;
reg [6:0] stripe_cnt;
reg [2:0] sub_h_cmp_g0;
reg [2:0] sub_h_cmp_g1;
reg [1:0] sub_h_cnt;
reg [2:0] sub_h_total_g0;
reg [2:0] sub_h_total_g1;
reg [2:0] sub_h_total_g10;
reg [2:0] sub_h_total_g11;
reg [1:0] sub_h_total_g2;
reg [2:0] sub_h_total_g3;
reg [2:0] sub_h_total_g4;
reg [2:0] sub_h_total_g5;
reg [2:0] sub_h_total_g6;
reg [2:0] sub_h_total_g7;
reg [2:0] sub_h_total_g8;
reg [2:0] sub_h_total_g9;
reg [13 -1:0] w_bias_d1;
reg [5:0] x_dilate;
reg [5:0] y_dilate;
wire [4:0] batch_cmp_w;
wire [4:0] batch_cnt_w;
wire [13 -1:0] c_bias_add;
wire c_bias_d1_reg_en;
wire c_bias_reg_en;
wire [13 -1:0] c_bias_w;
wire cbuf_reset;
wire [3:0] conv_x_stride_w;
wire [3:0] conv_y_stride_w;
wire dat_conv_req_dummy;
wire dat_dummy_l0_en;
wire dat_dummy_l1_en;
wire dat_dummy_l2_en;
wire dat_dummy_l3_en;
wire [15 -1:0] dat_entry_avl_add;
wire [15 -1:0] dat_entry_avl_sub;
wire [15 -1:0] dat_entry_avl_w;
wire [15 -1:0] dat_entry_end_inc;
wire [15 -1:0] dat_entry_end_inc_wrap;
wire [15 -1:0] dat_entry_end_w;
wire [15 -1:0] dat_entry_st_inc;
wire [15 -1:0] dat_entry_st_inc_wrap;
wire [15 -1:0] dat_entry_st_w;
wire mon_dat_entry_end_inc;
wire mon_dat_entry_st_inc;
wire dat_exec_valid;
wire dat_img_req_dummy;
wire dat_img_req_skip;
wire dat_l0_set;
wire dat_l0c0_dummy_w;
wire dat_l0c0_en;
wire dat_l0c1_dummy_w;
wire dat_l0c1_en;
wire dat_l1_set;
wire dat_l1c0_dummy_w;
wire dat_l1c0_en;
wire dat_l1c0_hi_en;
wire dat_l1c1_dummy_w;
wire dat_l1c1_en;
wire dat_l1c1_hi_en;
wire dat_l2_set;
wire dat_l2c0_dummy_w;
wire dat_l2c0_en;
wire dat_l2c1_dummy_w;
wire dat_l2c1_en;
wire dat_l3_set;
wire dat_l3c0_dummy_w;
wire dat_l3c0_en;
wire dat_l3c1_dummy_w;
wire dat_l3c1_en;
wire [512 -1:0] dat_out_bypass_data_w;
wire [64 -1:0] dat_out_bypass_mask_w;
wire dat_out_bypass_p0_vld_w;
wire [512 -1:0] dat_out_data;
wire [8:0] dat_out_flag_l0;
wire [8:0] dat_out_flag_w;
wire [64 -1:0] dat_out_mask;
wire dat_out_pvld_l0;
wire dat_out_pvld_w;
wire [512 -1:0] dat_out_wg_8b;
wire [512 -1:0] dat_out_wg_data;
wire [64 -1:0] dat_out_wg_mask;
wire [64 -1:0] dat_out_wg_mask_int8;
wire dat_pipe_local_valid_w;
wire dat_pipe_valid;
wire [512 -1:0] dat_pra_dat;
wire [255:0] dat_pra_dat_ch0;
wire [255:0] dat_pra_dat_ch1;
wire [255:0] dat_pra_dat_ch2;
wire [255:0] dat_pra_dat_ch3;
wire [13 -1:0] dat_req_addr_last;
wire [13:0] dat_req_addr_sum;
wire [13 -1:0] dat_req_addr_w;
wire [13 -1:0] dat_req_addr_wrap;
wire [13 -1:0] dat_req_base_d1;
wire mon_dat_req_addr_sum;
wire [4:0] dat_req_batch_index;
wire [7:0] dat_req_bytes;
wire dat_req_channel_end;
wire dat_req_dummy;
wire dat_req_exec_dummy;
wire dat_req_exec_pvld;
wire [1:0] dat_req_exec_sub_h;
wire [8:0] dat_req_flag_w;
wire dat_req_layer_end;
wire [7:0] dat_req_pipe_bytes;
wire dat_req_pipe_ch_end;
wire [1:0] dat_req_pipe_cur_sub_h;
wire dat_req_pipe_dummy;
wire [8:0] dat_req_pipe_flag;
wire [28:0] dat_req_pipe_pd;
wire dat_req_pipe_pvld;
wire dat_req_pipe_rls;
wire dat_req_pipe_sub_c;
wire [1:0] dat_req_pipe_sub_h;
wire [1:0] dat_req_pipe_sub_w;
wire dat_req_pipe_sub_w_st;
wire dat_req_skip;
wire dat_req_stripe_end;
wire dat_req_stripe_st;
wire dat_req_sub_c_w;
wire dat_req_sub_h_0_addr_en;
wire dat_req_sub_h_1_addr_en;
wire dat_req_sub_h_2_addr_en;
wire dat_req_sub_h_3_addr_en;
wire dat_req_sub_w_st_en;
wire [1:0] dat_req_sub_w_w;
wire dat_req_valid;
wire dat_rls;
wire [4:0] dat_rsp_batch_index;
wire [7:0] dat_rsp_bytes;
wire dat_rsp_ch_end;
wire dat_rsp_channel_end;
wire [512 -1:0] dat_rsp_conv;
wire [512 -1:0] dat_rsp_conv_8b;
wire [64 -1:0] dat_rsp_cur_h_e2_mask_8b;
wire [64 -1:0] dat_rsp_cur_h_e4_mask_8b;
wire [64 -1:0] dat_rsp_cur_h_mask_p1;
wire [31:0] dat_rsp_cur_h_mask_p2;
wire [31:0] dat_rsp_cur_h_mask_p3;
wire [1:0] dat_rsp_cur_sub_h;
wire [512 -1:0] dat_rsp_data_w;
wire dat_rsp_exec_dummy;
wire dat_rsp_exec_dummy_d0;
wire dat_rsp_exec_pvld;
wire dat_rsp_exec_pvld_d0;
wire [1:0] dat_rsp_exec_sub_h;
wire [1:0] dat_rsp_exec_sub_h_d0;
wire [8:0] dat_rsp_flag;
wire [512 -1:0] dat_rsp_img;
wire [512 -1:0] dat_rsp_img_8b;
wire dat_rsp_l0_block_end;
wire [8:0] dat_rsp_l0_flag;
wire dat_rsp_l0_pvld;
wire [512*2 -1:0] dat_rsp_l0_sft_in;
wire dat_rsp_l0_stripe_end;
wire dat_rsp_l0_sub_c;
wire [512 -1:0] dat_rsp_l0c0;
wire [512 -1:0] dat_rsp_l0c1;
wire dat_rsp_l1_block_end;
wire [8:0] dat_rsp_l1_flag;
wire dat_rsp_l1_pvld;
wire [512*2 -1:0] dat_rsp_l1_sft_in;
wire dat_rsp_l1_stripe_end;
wire dat_rsp_l1_sub_c;
wire [512 -1:0] dat_rsp_l1c0;
wire [512 -1:0] dat_rsp_l1c1;
wire dat_rsp_l2_block_end;
wire [8:0] dat_rsp_l2_flag;
wire dat_rsp_l2_pvld;
wire [512*2 -1:0] dat_rsp_l2_sft_in;
wire dat_rsp_l2_stripe_end;
wire dat_rsp_l2_sub_c;
wire [512 -1:0] dat_rsp_l2c0;
wire [512 -1:0] dat_rsp_l2c1;
wire dat_rsp_l3_block_end;
wire [8:0] dat_rsp_l3_flag;
wire dat_rsp_l3_pvld;
wire [512*2 -1:0] dat_rsp_l3_sft_in;
wire dat_rsp_l3_stripe_end;
wire dat_rsp_l3_sub_c;
wire [512 -1:0] dat_rsp_l3c0;
wire [512 -1:0] dat_rsp_l3c1;
wire dat_rsp_layer_end;
wire [64 -1:0] dat_rsp_mask_8b;
wire [64 -1:0] dat_rsp_mask_val_int8;
wire [64 -1:0] dat_rsp_mask_w;
wire [64 -1:0] dat_rsp_ori_mask;
wire dat_rsp_p0_vld_w;
wire dat_rsp_p1_vld_w;
wire [512 -1:0] dat_rsp_pad_value;
wire [26:0] dat_rsp_pd;
wire [26:0] dat_rsp_pd_d0;
wire [7:0] dat_rsp_pipe_bytes;
wire dat_rsp_pipe_ch_end;
wire [1:0] dat_rsp_pipe_cur_sub_h;
wire dat_rsp_pipe_dummy;
wire [8:0] dat_rsp_pipe_flag;
wire [28:0] dat_rsp_pipe_pd;
wire [28:0] dat_rsp_pipe_pd_d0;
wire dat_rsp_pipe_pvld;
wire dat_rsp_pipe_pvld_d0;
wire dat_rsp_pipe_rls;
wire dat_rsp_pipe_sub_c;
wire [1:0] dat_rsp_pipe_sub_h;
wire [1:0] dat_rsp_pipe_sub_w;
wire dat_rsp_pipe_sub_w_st;
wire dat_rsp_pra_en;
wire dat_rsp_pvld;
wire dat_rsp_pvld_d0;
wire dat_rsp_rls;
wire dat_rsp_stripe_end;
wire dat_rsp_stripe_st;
wire dat_rsp_sub_c;
wire [1:0] dat_rsp_sub_h;
wire [1:0] dat_rsp_sub_w;
wire [512 -1:0] dat_rsp_wg;
wire [255:0] dat_rsp_wg_ch0;
wire [255:0] dat_rsp_wg_ch1;
wire [255:0] dat_rsp_wg_ch2;
wire [255:0] dat_rsp_wg_ch3;
wire [512 -1:0] dat_rsp_wg_lb;
wire [512 -1:0] dat_rsp_wg_lt;
wire [512 -1:0] dat_rsp_wg_rb;
wire [512 -1:0] dat_rsp_wg_rt;
wire dat_rsp_wg_sel_8b_hi;
wire dat_rsp_wg_sel_8b_lo;
wire dat_rsp_wg_sel_lb;
wire dat_rsp_wg_sel_lt;
wire dat_rsp_wg_sel_rb;
wire dat_rsp_wg_sel_rt;
wire [13:0] dat_slice_avl_add;
wire [13:0] dat_slice_avl_sub;
wire [13:0] dat_slice_avl_w;
wire [2303:0] dat_wg;
wire [255:0] dat_wg_8b_ch0;
wire [255:0] dat_wg_8b_ch1;
wire [255:0] dat_wg_8b_ch2;
wire [255:0] dat_wg_8b_ch3;
wire [255:0] dat_wg_8b_ch4;
wire [255:0] dat_wg_8b_ch5;
wire [255:0] dat_wg_8b_ch6;
wire [255:0] dat_wg_8b_ch7;
wire dat_wg_adv;
wire dat_wg_req_dummy;
wire dat_wg_req_skip;
wire [4:0] data_bank_w;
wire [5:0] data_batch_w;
wire [10:0] datain_c_cnt_inc;
wire datain_c_cnt_reg_en;
wire [10:0] datain_c_cnt_w;
wire [10:0] datain_channel_cmp_w;
wire [13:0] datain_h_cnt_inc;
wire datain_h_cnt_reg_en;
wire [13:0] datain_h_cnt_st;
wire [13:0] datain_h_cnt_w;
wire [13:0] datain_h_cur;
wire datain_h_ori_reg_en;
wire [12:0] datain_height_cmp_w;
wire [13:0] datain_w_cnt_inc;
wire datain_w_cnt_reg_en;
wire [13:0] datain_w_cnt_st;
wire [13:0] datain_w_cnt_w;
wire [13:0] datain_w_cur;
wire datain_w_ori_reg_en;
wire [12:0] datain_width_cmp_w;
wire [13:0] datain_width_w;
wire [2:0] dataout_w_add;
wire [12:0] dataout_w_cnt_inc;
wire dataout_w_cnt_reg_en;
wire [12:0] dataout_w_cnt_w;
wire [12:0] dataout_w_init;
wire dataout_w_ori_reg_en;
wire [12:0] dataout_width_cmp_w;
wire [512 -1:0] dbg_csc_dat;
//: for(my $i=0; $i<64 ; $i++){
//: print qq(
//: wire [8 -1:0] dbg_csc_dat_${i}; )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

wire [8 -1:0] dbg_csc_dat_0; 
wire [8 -1:0] dbg_csc_dat_1; 
wire [8 -1:0] dbg_csc_dat_2; 
wire [8 -1:0] dbg_csc_dat_3; 
wire [8 -1:0] dbg_csc_dat_4; 
wire [8 -1:0] dbg_csc_dat_5; 
wire [8 -1:0] dbg_csc_dat_6; 
wire [8 -1:0] dbg_csc_dat_7; 
wire [8 -1:0] dbg_csc_dat_8; 
wire [8 -1:0] dbg_csc_dat_9; 
wire [8 -1:0] dbg_csc_dat_10; 
wire [8 -1:0] dbg_csc_dat_11; 
wire [8 -1:0] dbg_csc_dat_12; 
wire [8 -1:0] dbg_csc_dat_13; 
wire [8 -1:0] dbg_csc_dat_14; 
wire [8 -1:0] dbg_csc_dat_15; 
wire [8 -1:0] dbg_csc_dat_16; 
wire [8 -1:0] dbg_csc_dat_17; 
wire [8 -1:0] dbg_csc_dat_18; 
wire [8 -1:0] dbg_csc_dat_19; 
wire [8 -1:0] dbg_csc_dat_20; 
wire [8 -1:0] dbg_csc_dat_21; 
wire [8 -1:0] dbg_csc_dat_22; 
wire [8 -1:0] dbg_csc_dat_23; 
wire [8 -1:0] dbg_csc_dat_24; 
wire [8 -1:0] dbg_csc_dat_25; 
wire [8 -1:0] dbg_csc_dat_26; 
wire [8 -1:0] dbg_csc_dat_27; 
wire [8 -1:0] dbg_csc_dat_28; 
wire [8 -1:0] dbg_csc_dat_29; 
wire [8 -1:0] dbg_csc_dat_30; 
wire [8 -1:0] dbg_csc_dat_31; 
wire [8 -1:0] dbg_csc_dat_32; 
wire [8 -1:0] dbg_csc_dat_33; 
wire [8 -1:0] dbg_csc_dat_34; 
wire [8 -1:0] dbg_csc_dat_35; 
wire [8 -1:0] dbg_csc_dat_36; 
wire [8 -1:0] dbg_csc_dat_37; 
wire [8 -1:0] dbg_csc_dat_38; 
wire [8 -1:0] dbg_csc_dat_39; 
wire [8 -1:0] dbg_csc_dat_40; 
wire [8 -1:0] dbg_csc_dat_41; 
wire [8 -1:0] dbg_csc_dat_42; 
wire [8 -1:0] dbg_csc_dat_43; 
wire [8 -1:0] dbg_csc_dat_44; 
wire [8 -1:0] dbg_csc_dat_45; 
wire [8 -1:0] dbg_csc_dat_46; 
wire [8 -1:0] dbg_csc_dat_47; 
wire [8 -1:0] dbg_csc_dat_48; 
wire [8 -1:0] dbg_csc_dat_49; 
wire [8 -1:0] dbg_csc_dat_50; 
wire [8 -1:0] dbg_csc_dat_51; 
wire [8 -1:0] dbg_csc_dat_52; 
wire [8 -1:0] dbg_csc_dat_53; 
wire [8 -1:0] dbg_csc_dat_54; 
wire [8 -1:0] dbg_csc_dat_55; 
wire [8 -1:0] dbg_csc_dat_56; 
wire [8 -1:0] dbg_csc_dat_57; 
wire [8 -1:0] dbg_csc_dat_58; 
wire [8 -1:0] dbg_csc_dat_59; 
wire [8 -1:0] dbg_csc_dat_60; 
wire [8 -1:0] dbg_csc_dat_61; 
wire [8 -1:0] dbg_csc_dat_62; 
wire [8 -1:0] dbg_csc_dat_63; 
//| eperl: generated_end (DO NOT EDIT ABOVE)
wire dl_block_end;
wire dl_channel_end;
wire [6:0] dl_channel_size;
wire [1:0] dl_cur_sub_h;
wire dl_dat_release;
wire dl_group_end;
wire [4:0] dl_h_offset;
wire [9:0] dl_h_offset_ext;
wire [30:0] dl_in_pd;
wire [30:0] dl_in_pd_d0;
wire dl_in_pvld;
wire dl_in_pvld_d0;
wire dl_layer_end;
wire [30:0] dl_pd;
wire [30:0] dl_pd_d0;
wire dl_pvld;
wire dl_pvld_d0;
wire [6:0] dl_stripe_length;
wire [4:0] dl_w_offset;
wire [9:0] dl_w_offset_ext;
wire [15 -1:0] entries_batch_w;
wire [15 -1:0] entries_single_w;
wire [15 -1:0] entries_w;
wire [13 -1:0] h_bias_0_stride_w;
wire [13 -1:0] h_bias_0_w;
wire [13 -1:0] h_bias_1_stride_w;
wire [13 -1:0] h_bias_1_w;
wire [13 -1:0] h_bias_2_w;
wire [13 -1:0] h_bias_3_w;
wire [13 -1:0] h_bias_d1;
wire [1:0] h_bias_reg_en;
wire [13:0] h_offset_slice_w;
wire is_batch_end;
wire is_conv;
wire is_dat_entry_end_wrap;
wire is_dat_entry_st_wrap;
wire is_dat_req_addr_wrap;
wire is_img;
wire is_last_channel;
wire is_pixel;
wire is_running_first;
wire is_sg_done;
wire is_sg_idle;
wire is_sg_running;
wire is_stripe_end;
wire is_stripe_equal;
wire is_sub_h_end;
wire is_w_end;
wire is_w_end_ahead;
wire is_winograd;
wire layer_st;
wire mon_batch_cnt_w;
wire mon_c_bias_w;
wire mon_dat_entry_avl_w;
wire mon_dat_entry_end_inc_wrap;
wire mon_dat_entry_st_inc_wrap;
wire [3:0] mon_dat_out_pra_vld;
wire [1:0] mon_dat_req_addr_wrap;
wire [512 -1:0] mon_dat_rsp_l0_sft;
wire [512 -1:0] mon_dat_rsp_l1_sft;
wire [512 -1:0] mon_dat_rsp_l2_sft;
wire [512 -1:0] mon_dat_rsp_l3_sft;
wire [3:0] mon_dat_rsp_pra_rdy;
wire mon_dat_slice_avl_w;
wire mon_data_bank_w;
wire mon_datain_c_cnt_inc;
wire mon_datain_h_cnt_inc;
wire mon_datain_h_cur;
wire mon_datain_w_cnt_inc;
wire mon_datain_w_cur;
wire mon_dataout_w_cnt_inc;
wire [5:0] mon_entries_batch_w;
wire mon_entries_single_w;
wire mon_entries_w;
wire [5:0] mon_h_bias_0_stride_w;
wire [13 -1:0] mon_h_bias_0_w;
wire [12:0] mon_h_bias_1_stride_w;
wire [4:0] mon_h_bias_1_w;
wire [4:0] mon_h_bias_2_w;
wire [1:0] mon_h_bias_3_w;
wire mon_h_bias_d1;
wire mon_pixel_w_cnt_w;
wire [1:0] mon_pixel_x_init_w;
wire mon_rls_slices_w;
wire mon_rsp_sft_cnt_l0_w;
wire mon_rsp_sft_cnt_l1_w;
wire mon_rsp_sft_cnt_l2_w;
wire mon_rsp_sft_cnt_l3_w;
wire [13:0] mon_slice_entries_w;
wire [1:0] mon_slice_left_w;
wire mon_stripe_cnt_inc;
wire [2:0] mon_sub_h_total_w;
wire pixel_ch_ori_reg_en;
wire [11:0] pixel_ch_stride_w;
wire pixel_force_clr;
wire pixel_force_fetch;
wire pixel_w_cnt_reg_en;
wire [15:0] pixel_w_cnt_w;
wire [14:0] pixel_w_cur;
wire pixel_w_ori_reg_en;
wire [7:0] pixel_x_add_w;
wire [6:0] pixel_x_byte_stride_w;
wire [6:0] pixel_x_cnt_add;
wire [6:0] pixel_x_init_offset_w;
wire [5:0] pixel_x_init_w;
wire [5:0] pixel_x_stride_w;
wire [1:0] pra_precision_0;
wire [1:0] pra_precision_1;
wire [1:0] pra_precision_2;
wire [1:0] pra_precision_3;
wire [1:0] pra_truncate_0;
wire [1:0] pra_truncate_1;
wire [1:0] pra_truncate_2;
wire [1:0] pra_truncate_3;
wire [1:0] pra_truncate_w;
wire reuse_rls;
wire [13:0] rls_slices_w;
wire rsp_sft_cnt_l0_en;
wire [7:0] rsp_sft_cnt_l0_inc;
wire rsp_sft_cnt_l0_ori_en;
wire [7:0] rsp_sft_cnt_l0_sub;
wire [7:0] rsp_sft_cnt_l0_w;
wire rsp_sft_cnt_l1_en;
wire [7:0] rsp_sft_cnt_l1_inc;
wire rsp_sft_cnt_l1_ori_en;
wire [7:0] rsp_sft_cnt_l1_sub;
wire [7:0] rsp_sft_cnt_l1_w;
wire rsp_sft_cnt_l2_en;
wire [7:0] rsp_sft_cnt_l2_inc;
wire rsp_sft_cnt_l2_ori_en;
wire [7:0] rsp_sft_cnt_l2_sub;
wire [7:0] rsp_sft_cnt_l2_w;
wire rsp_sft_cnt_l3_en;
wire [7:0] rsp_sft_cnt_l3_inc;
wire rsp_sft_cnt_l3_ori_en;
wire [7:0] rsp_sft_cnt_l3_sub;
wire [7:0] rsp_sft_cnt_l3_w;
wire rsp_sft_l1_sel_1;
wire rsp_sft_l1_sel_2;
wire rsp_sft_l1_sel_3;
wire rsp_sft_l2_sel_1;
wire rsp_sft_l2_sel_2;
wire rsp_sft_l2_sel_3;
wire rsp_sft_l3_sel_1;
wire rsp_sft_l3_sel_2;
wire rsp_sft_l3_sel_3;
wire sc2buf_dat_rd_en_w;
wire [15 -1:0] sc2cdma_dat_entries_w;
wire [13:0] sc2cdma_dat_slices_w;
wire [8:0] sc2mac_dat_pd_w;
wire slcg_wg_en_w;
wire [15 -1:0] slice_entries_w;
wire [13:0] slice_left_w;
wire [13:0] slices_oprand;
wire [6:0] stripe_cnt_inc;
wire stripe_cnt_reg_en;
wire [6:0] stripe_cnt_w;
wire [2:0] sub_h_cmp_w;
wire [2:0] sub_h_cnt_inc;
wire sub_h_cnt_reg_en;
wire [1:0] sub_h_cnt_w;
wire [2:0] sub_h_total_w;
wire sub_rls;
wire [14:0] w_bias_int8;
wire w_bias_reg_en;
wire [13:0] w_bias_w;
wire [5:0] x_dilate_w;
wire [5:0] y_dilate_w;
/////////////////////////////////////////////////////////////////////////////////////////////
// Pipeline of Weight loader, for both compressed weight and uncompressed weight
//
// input_package
// |
// data request
// |
// conv_buffer
// |
// feature data---> data relase
// | |
// REG PRA
// | |
// REGISTER
// |
// MAC
//
/////////////////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////
///// status from sequence generator                     /////
//////////////////////////////////////////////////////////////
assign is_sg_idle = (sc_state == 0 );
assign is_sg_running = (sc_state == 2 );
assign is_sg_done = (sc_state == 3 );
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"is_sg_running\" -q is_sg_running_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       is_sg_running_d1 <= 1'b0;
   end else begin
       is_sg_running_d1 <= is_sg_running;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// input signals from registers                       /////
//////////////////////////////////////////////////////////////
assign layer_st = reg2dp_op_en & is_sg_idle;
assign is_pixel = (reg2dp_datain_format == 1'h1 );
assign is_winograd = 1'b0;
assign is_conv = (reg2dp_conv_mode == 1'h0 );
assign is_img = is_conv & is_pixel;
assign {mon_data_bank_w, data_bank_w} = reg2dp_data_bank + 1'b1;
assign data_batch_w = 6'b1;
assign batch_cmp_w = 5'b0;
//assign is_int8 = (reg2dp_proc_precision == 2'h0 );
//assign is_fp16 = (reg2dp_proc_precision == 2'h2 );
assign datain_width_w = is_winograd ? ({2'b0, reg2dp_datain_width_ext[12:2]} + 1'b1) : reg2dp_datain_width_ext + 1'b1;
assign datain_width_cmp_w = reg2dp_datain_width_ext;
assign datain_height_cmp_w = reg2dp_datain_height_ext;
assign datain_channel_cmp_w = is_winograd ? reg2dp_weight_channel_ext[12:2] : {{6 -2{1'b0}}, reg2dp_weight_channel_ext[12:6]};
//y_ex=0,sub_h_total=1;y_ex=1,sub_h_total=2; y_ext=2,sub_h_total=4; non_image, sub_h_total=1;
//sub_h_total means how many h lines are used in post-extention
assign {sub_h_total_w, mon_sub_h_total_w} = is_img ? (6'h9 << reg2dp_y_extension) : 6'h8;
assign sub_h_cmp_w = is_img ? sub_h_total_w : is_winograd ? 3'h2 : 3'h1;
assign dataout_w_init[12:0] = sub_h_cmp_w - 1'b1;
assign conv_x_stride_w = (is_winograd) ? 4'b1 : reg2dp_conv_x_stride_ext + 1'b1;
assign pixel_x_stride_w = (reg2dp_datain_channel_ext[1:0] == 2'h3) ? {conv_x_stride_w, 2'b0} : //*4, after pre_extension
                          (reg2dp_datain_channel_ext[1:0] == 2'h2) ? ({conv_x_stride_w, 1'b0} + conv_x_stride_w) : //*3
                          {2'b0, conv_x_stride_w}; //*1
//: my $kk=6;
//: if ($kk=6) {
//: print qq (
//: assign {mon_pixel_x_init_w,pixel_x_init_w} = (reg2dp_y_extension == 2'h2) ? ({pixel_x_stride_w, 1'b0} + pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]) :
//: (reg2dp_y_extension == 2'h1) ? (pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]):
//: (reg2dp_weight_channel_ext >= 7'h40) ? {6{1'b1}}: //cut by atomC
//: {reg2dp_weight_channel_ext[6 -1:0]};
//: )
//: }
//: else {
//: print qq(
//: assign {mon_pixel_x_init_w,pixel_x_init_w} = (reg2dp_y_extension == 2'h2) ? ({pixel_x_stride_w, 1'b0} + pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]) :
//: (reg2dp_y_extension == 2'h1) ? (pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]):
//: (reg2dp_weight_channel_ext >= 7'h40) ? {6{1'b1}}: //cut by atomC
//: {{6-6{1'b0}},reg2dp_weight_channel_ext[6 -1:0]};
//: )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

assign {mon_pixel_x_init_w,pixel_x_init_w} = (reg2dp_y_extension == 2'h2) ? ({pixel_x_stride_w, 1'b0} + pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]) :
(reg2dp_y_extension == 2'h1) ? (pixel_x_stride_w + reg2dp_weight_channel_ext[5:0]):
(reg2dp_weight_channel_ext >= 7'h40) ? {6{1'b1}}: //cut by atomC
{reg2dp_weight_channel_ext[6 -1:0]};

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign pixel_x_init_offset_w = (reg2dp_weight_channel_ext[6 -1:0] + 1'b1);
assign pixel_x_add_w = (reg2dp_y_extension == 2'h2) ? {pixel_x_stride_w, 2'b0} : //*4, after post_extension
                       (reg2dp_y_extension == 2'h1) ? {1'b0, pixel_x_stride_w, 1'b0} : //*2
                       {2'b0, pixel_x_stride_w};
assign pixel_x_byte_stride_w = {1'b0, pixel_x_stride_w};
//: my $kk=5;
//: if($kk=5) {
//: print qq(
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_1
//: assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_2
//: assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_4
//: assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +2{1'b0}}}; //stick to 4*atomK  no matter which config.  
//: `endif
//: )
//: }
//: else {
//: print qq(
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_1
//: assign pixel_ch_stride_w = {{5-5{1'b0}},pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_2
//: assign pixel_ch_stride_w = {{5-5{1'b0}},pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  
//: `endif
//: `ifdef CC_ATOMC_DIV_ATOMK_EQUAL_4
//: assign pixel_ch_stride_w = {{5-5{1'b0}},pixel_x_stride_w, {5 +2{1'b0}}}; //stick to 4*atomK  no matter which config.  
//: `endif
//: )
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)

assign pixel_ch_stride_w = {pixel_x_stride_w, {5 +1{1'b0}}}; //stick to 2*atomK  no matter which config.  


//| eperl: generated_end (DO NOT EDIT ABOVE)
assign conv_y_stride_w = (is_winograd) ? 4'b1 : reg2dp_conv_y_stride_ext + 1'b1;
assign x_dilate_w = (is_winograd | is_img) ? 6'b1 : reg2dp_x_dilation_ext + 1'b1;
assign y_dilate_w = (is_winograd | is_img) ? 6'b1 : reg2dp_y_dilation_ext + 1'b1;
//reg2dp_entries means entry per slice
assign {mon_entries_single_w,entries_single_w} = (reg2dp_entries + 1'b1);
assign {mon_entries_batch_w,entries_batch_w} = entries_single_w * data_batch_w;
assign {mon_entries_w,entries_w} = (is_winograd) ? ({reg2dp_entries[12:0], 2'b0} + 3'h4) : entries_single_w;
assign h_offset_slice_w[11:0] = data_batch_w * y_dilate_w;
assign h_offset_slice_w[13:12] = 2'b0;
assign {mon_h_bias_0_stride_w,h_bias_0_stride_w} = entries * data_batch;
assign {mon_h_bias_1_stride_w,h_bias_1_stride_w} = entries * h_offset_slice;
assign {mon_rls_slices_w,rls_slices_w} = reg2dp_rls_slices + 1'b1;
assign {mon_slice_left_w,slice_left_w} = reg2dp_skip_data_rls ? (reg2dp_datain_height_ext + 1'b1) : reg2dp_datain_height_ext - reg2dp_rls_slices;
assign slices_oprand = layer_st_d1 ? rls_slices : slice_left;
assign {mon_slice_entries_w,slice_entries_w} = entries_batch * slices_oprand;
assign dataout_width_cmp_w = reg2dp_dataout_width;
assign pra_truncate_w = (reg2dp_pra_truncate == 2'h3) ? 2'h2 : reg2dp_pra_truncate;
//: my $kk=15;
//: my $jj=13;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"layer_st\" -q layer_st_d1");
//: &eperl::flop("-nodeclare   -rval \"{22{1'b0}}\"  -en \"layer_st\" -d \"{22{is_winograd}}\" -q is_winograd_d1");
//: &eperl::flop("-nodeclare   -rval \"{34{1'b0}}\"  -en \"layer_st\" -d \"{34{is_img}}\" -q is_img_d1");
//: &eperl::flop("-nodeclare   -rval \"{5{1'b0}}\"  -en \"layer_st\" -d \"data_bank_w\" -q data_bank");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"datain_width_w\" -q datain_width");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"layer_st\" -d \"datain_width_cmp_w\" -q datain_width_cmp");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"layer_st\" -d \"datain_height_cmp_w\" -q datain_height_cmp");
//: &eperl::flop("-nodeclare   -rval \"{11{1'b0}}\"  -en \"layer_st\" -d \"datain_channel_cmp_w\" -q datain_channel_cmp");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g0");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g1");
//: &eperl::flop("-nodeclare   -rval \"2'h1\"  -en \"layer_st\" -d \"sub_h_total_w[2:1]\" -q sub_h_total_g2");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g3");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g4");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g5");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g6");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g7");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g8");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g9");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g10");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_total_w\" -q sub_h_total_g11");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_cmp_w\" -q sub_h_cmp_g0");
//: &eperl::flop("-nodeclare   -rval \"3'h1\"  -en \"layer_st\" -d \"sub_h_cmp_w\" -q sub_h_cmp_g1");
//: &eperl::flop("-nodeclare   -rval \"{4{1'b0}}\"  -en \"layer_st\" -d \"conv_x_stride_w\" -q conv_x_stride");
//: &eperl::flop("-nodeclare   -rval \"{4{1'b0}}\"  -en \"layer_st\" -d \"conv_y_stride_w\" -q conv_y_stride");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"layer_st\" -d \"pixel_x_stride_w[0]\" -q pixel_x_stride_odd");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"data_batch_w\" -q data_batch");
//: &eperl::flop("-nodeclare   -rval \"{5{1'b0}}\"  -en \"layer_st\" -d \"batch_cmp_w\" -q batch_cmp");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_init_w\" -q pixel_x_init");
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_init_offset_w\" -q pixel_x_init_offset");
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_add_w[6:0]\" -q pixel_x_add");
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"layer_st\" -d \"pixel_x_byte_stride_w\" -q pixel_x_byte_stride");
//: &eperl::flop("-nodeclare   -rval \"{12{1'b0}}\"  -en \"layer_st\" -d \"pixel_ch_stride_w\" -q pixel_ch_stride");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"x_dilate_w\" -q x_dilate");
//: &eperl::flop("-nodeclare   -rval \"{6{1'b0}}\"  -en \"layer_st\" -d \"y_dilate_w\" -q y_dilate");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"layer_st\" -d \"reg2dp_pad_value\" -q pad_value");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st\" -d \"entries_w\" -q entries");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st\" -d \"entries_batch_w\" -q entries_batch");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st\" -d \"{1'h0,reg2dp_entries}\" -q entries_cmp");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"h_offset_slice_w\" -q h_offset_slice");
//: &eperl::flop("-nodeclare   -rval \"{12{1'b0}}\"  -en \"layer_st_d1\" -d \"h_bias_0_stride_w\" -q h_bias_0_stride");
//: &eperl::flop("-nodeclare   -rval \"{12{1'b0}}\"  -en \"layer_st_d1\" -d \"h_bias_1_stride_w\" -q h_bias_1_stride");
//: &eperl::flop("-nodeclare   -rval \"{${jj}{1'b0}}\"  -en \"layer_st_d1\" -d \"entries[${jj}-1:0]\" -q h_bias_2_stride");
//: &eperl::flop("-nodeclare   -rval \"{${jj}{1'b0}}\"  -en \"layer_st_d1\" -d \"entries[${jj}-1:0]\" -q h_bias_3_stride");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"rls_slices_w\" -q rls_slices");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"layer_st_d1\" -d \"slice_entries_w\" -q rls_entries");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"layer_st\" -d \"slice_left_w[13:0]\" -q slice_left");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"is_sg_done\" -d \"slice_left\" -q last_slices");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"is_sg_done\" -d \"slice_entries_w\" -q last_entries");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"layer_st\" -d \"dataout_width_cmp_w\" -q dataout_width_cmp");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"layer_st\" -d \"{4{pra_truncate_w}}\" -q pra_truncate");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"layer_st\" -d \"{4{reg2dp_proc_precision}}\" -q pra_precision");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       layer_st_d1 <= 1'b0;
   end else begin
       layer_st_d1 <= layer_st;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       is_winograd_d1 <= {22{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           is_winograd_d1 <= {22{is_winograd}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           is_winograd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       is_img_d1 <= {34{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           is_img_d1 <= {34{is_img}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           is_img_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       data_bank <= {5{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           data_bank <= data_bank_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           data_bank <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_width <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_width <= datain_width_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_width <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_width_cmp <= {13{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_width_cmp <= datain_width_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_width_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_height_cmp <= {13{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_height_cmp <= datain_height_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_height_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_channel_cmp <= {11{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           datain_channel_cmp <= datain_channel_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           datain_channel_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g0 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g0 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g0 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g1 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g1 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g2 <= 2'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g2 <= sub_h_total_w[2:1];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g3 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g3 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g4 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g4 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g4 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g5 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g5 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g5 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g6 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g6 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g6 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g7 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g7 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g7 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g8 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g8 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g8 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g9 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g9 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g9 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g10 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g10 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g10 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_total_g11 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_total_g11 <= sub_h_total_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_total_g11 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_cmp_g0 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_cmp_g0 <= sub_h_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_cmp_g0 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_cmp_g1 <= 3'h1;
   end else begin
       if ((layer_st) == 1'b1) begin
           sub_h_cmp_g1 <= sub_h_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           sub_h_cmp_g1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       conv_x_stride <= {4{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           conv_x_stride <= conv_x_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           conv_x_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       conv_y_stride <= {4{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           conv_y_stride <= conv_y_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           conv_y_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_stride_odd <= 1'b0;
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_stride_odd <= pixel_x_stride_w[0];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_stride_odd <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       data_batch <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           data_batch <= data_batch_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           data_batch <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       batch_cmp <= {5{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           batch_cmp <= batch_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           batch_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_init <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_init <= pixel_x_init_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_init <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_init_offset <= {7{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_init_offset <= pixel_x_init_offset_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_init_offset <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_add <= {7{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_add <= pixel_x_add_w[6:0];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_add <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_x_byte_stride <= {7{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_x_byte_stride <= pixel_x_byte_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_x_byte_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_ch_stride <= {12{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pixel_ch_stride <= pixel_ch_stride_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pixel_ch_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       x_dilate <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           x_dilate <= x_dilate_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           x_dilate <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       y_dilate <= {6{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           y_dilate <= y_dilate_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           y_dilate <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pad_value <= {16{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pad_value <= reg2dp_pad_value;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pad_value <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       entries <= {15{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           entries <= entries_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           entries <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       entries_batch <= {15{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           entries_batch <= entries_batch_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           entries_batch <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       entries_cmp <= {15{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           entries_cmp <= {1'h0,reg2dp_entries};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           entries_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_offset_slice <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           h_offset_slice <= h_offset_slice_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           h_offset_slice <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_0_stride <= {12{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_0_stride <= h_bias_0_stride_w;
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_0_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_1_stride <= {12{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_1_stride <= h_bias_1_stride_w;
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_1_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_2_stride <= {13{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_2_stride <= entries[13-1:0];
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_2_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_3_stride <= {13{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           h_bias_3_stride <= entries[13-1:0];
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           h_bias_3_stride <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rls_slices <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           rls_slices <= rls_slices_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           rls_slices <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rls_entries <= {15{1'b0}};
   end else begin
       if ((layer_st_d1) == 1'b1) begin
           rls_entries <= slice_entries_w;
       // VCS coverage off
       end else if ((layer_st_d1) == 1'b0) begin
       end else begin
           rls_entries <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slice_left <= {14{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           slice_left <= slice_left_w[13:0];
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           slice_left <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       last_slices <= {14{1'b0}};
   end else begin
       if ((is_sg_done) == 1'b1) begin
           last_slices <= slice_left;
       // VCS coverage off
       end else if ((is_sg_done) == 1'b0) begin
       end else begin
           last_slices <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       last_entries <= {15{1'b0}};
   end else begin
       if ((is_sg_done) == 1'b1) begin
           last_entries <= slice_entries_w;
       // VCS coverage off
       end else if ((is_sg_done) == 1'b0) begin
       end else begin
           last_entries <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dataout_width_cmp <= {13{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           dataout_width_cmp <= dataout_width_cmp_w;
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           dataout_width_cmp <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pra_truncate <= {8{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pra_truncate <= {4{pra_truncate_w}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pra_truncate <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pra_precision <= {8{1'b0}};
   end else begin
       if ((layer_st) == 1'b1) begin
           pra_precision <= {4{reg2dp_proc_precision}};
       // VCS coverage off
       end else if ((layer_st) == 1'b0) begin
       end else begin
           pra_precision <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////////////////////////////////////////////////////
// SLCG control signal //
////////////////////////////////////////////////////////////////////////
assign slcg_wg_en_w = reg2dp_op_en & is_winograd;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"slcg_wg_en_w\" -q slcg_wg_en_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"slcg_wg_en_d1\" -q slcg_wg_en_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"slcg_wg_en_d2\" -q slcg_wg_en_d3");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slcg_wg_en_d1 <= 1'b0;
   end else begin
       slcg_wg_en_d1 <= slcg_wg_en_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slcg_wg_en_d2 <= 1'b0;
   end else begin
       slcg_wg_en_d2 <= slcg_wg_en_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       slcg_wg_en_d3 <= 1'b0;
   end else begin
       slcg_wg_en_d3 <= slcg_wg_en_d2;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign slcg_wg_en = slcg_wg_en_d3;
//////////////////////////////////////////////////////////////
///// cbuf status management                             /////
//////////////////////////////////////////////////////////////
//================ Non-SLCG clock domain ================//
assign cbuf_reset = sc2cdma_dat_pending_req;
assign is_running_first = is_sg_running & ~is_sg_running_d1;
//////////////////////////////////// calculate how many avaliable dat slices in cbuf////////////////////////////////////
assign dat_slice_avl_add = cdma2sc_dat_updt ? cdma2sc_dat_slices : 14'b0;
assign dat_slice_avl_sub = dat_rls ? sc2cdma_dat_slices_w : 14'b0;
assign {mon_dat_slice_avl_w, dat_slice_avl_w} = (cbuf_reset) ? 14'b0 : dat_slice_avl + dat_slice_avl_add - dat_slice_avl_sub;
//////////////////////////////////// calculate how many avaliable dat entries in cbuf////////////////////////////////////
assign dat_entry_avl_add = cdma2sc_dat_updt ? cdma2sc_dat_entries :{15{1'b0}};
assign dat_entry_avl_sub = dat_rls ? sc2cdma_dat_entries_w : {15{1'b0}};
assign {mon_dat_entry_avl_w,dat_entry_avl_w} = (cbuf_reset) ? {15{1'b0}} : dat_entry_avl + dat_entry_avl_add - dat_entry_avl_sub;
//////////////////////////////////// calculate avilable data entries start offset in cbuf banks ////////////////////////////////////
// data_bank is the highest bank for storing data
assign {mon_dat_entry_st_inc,dat_entry_st_inc} = dat_entry_st + dat_entry_avl_sub;
assign {mon_dat_entry_st_inc_wrap, dat_entry_st_inc_wrap} = dat_entry_st_inc - {data_bank, {9{1'b0}} };
assign is_dat_entry_st_wrap = (dat_entry_st_inc >= {1'b0, data_bank, {9{1'b0}} });
assign dat_entry_st_w = (cbuf_reset) ? {15{1'b0}} : is_dat_entry_st_wrap ? dat_entry_st_inc_wrap : dat_entry_st_inc[15 -1:0];
//////////////////////////////////// calculate avilable data entries end offset in cbuf banks////////////////////////////////////
assign {mon_dat_entry_end_inc,dat_entry_end_inc} = dat_entry_end + dat_entry_avl_add;
assign {mon_dat_entry_end_inc_wrap,dat_entry_end_inc_wrap} = dat_entry_end_inc - {data_bank, {9{1'b0}} };
assign is_dat_entry_end_wrap = (dat_entry_end_inc >= {1'b0, data_bank, {9{1'b0}} });
assign dat_entry_end_w = (cbuf_reset) ? {15{1'b0}} : is_dat_entry_end_wrap ? dat_entry_end_inc_wrap : dat_entry_end_inc[15 -1:0];
//////////////////////////////////// registers and assertions ////////////////////////////////////
//: my $kk= 15;
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{14{1'b0}}\"  -en \"cdma2sc_dat_updt | dat_rls | cbuf_reset\" -d \"dat_slice_avl_w\" -q dat_slice_avl");
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{${kk}{1'b0}}\"  -en \"cdma2sc_dat_updt | dat_rls | cbuf_reset\" -d \"dat_entry_avl_w\" -q dat_entry_avl");
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{${kk}{1'b0}}\"  -en \"cbuf_reset | dat_rls\" -d \"dat_entry_st_w\" -q dat_entry_st");
//: &eperl::flop("-nodeclare -clk nvdla_core_ng_clk  -rval \"{${kk}{1'b0}}\"  -en \"cbuf_reset | cdma2sc_dat_updt\" -d \"dat_entry_end_w\" -q dat_entry_end");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_ng_clk) begin
   if (!nvdla_core_rstn) begin
       dat_slice_avl <= {14{1'b0}};
   end else begin
       if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b1) begin
           dat_slice_avl <= dat_slice_avl_w;
       // VCS coverage off
       end else if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b0) begin
       end else begin
           dat_slice_avl <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_ng_clk) begin
   if (!nvdla_core_rstn) begin
       dat_entry_avl <= {15{1'b0}};
   end else begin
       if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b1) begin
           dat_entry_avl <= dat_entry_avl_w;
       // VCS coverage off
       end else if ((cdma2sc_dat_updt | dat_rls | cbuf_reset) == 1'b0) begin
       end else begin
           dat_entry_avl <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_ng_clk) begin
   if (!nvdla_core_rstn) begin
       dat_entry_st <= {15{1'b0}};
   end else begin
       if ((cbuf_reset | dat_rls) == 1'b1) begin
           dat_entry_st <= dat_entry_st_w;
       // VCS coverage off
       end else if ((cbuf_reset | dat_rls) == 1'b0) begin
       end else begin
           dat_entry_st <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_ng_clk) begin
   if (!nvdla_core_rstn) begin
       dat_entry_end <= {15{1'b0}};
   end else begin
       if ((cbuf_reset | cdma2sc_dat_updt) == 1'b1) begin
           dat_entry_end <= dat_entry_end_w;
       // VCS coverage off
       end else if ((cbuf_reset | cdma2sc_dat_updt) == 1'b0) begin
       end else begin
           dat_entry_end <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//================ Non-SLCG clock domain end ================//
//////////////////////////////////////////////////////////////
///// cbuf status update                                 /////
//////////////////////////////////////////////////////////////
assign sub_rls = (dat_rsp_pvld & dat_rsp_rls);
assign reuse_rls = sg2dl_reuse_rls;
assign dat_rls = (reuse_rls & (|last_slices)) | (sub_rls & (|rls_slices));
assign sc2cdma_dat_slices_w = sub_rls ? rls_slices : last_slices;
assign sc2cdma_dat_entries_w = sub_rls ? rls_entries : last_entries;
//: my $kk=15;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_rls\" -q sc2cdma_dat_updt");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"dat_rls\" -d \"sc2cdma_dat_slices_w[13:0]\" -q sc2cdma_dat_slices");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dat_rls\" -d \"sc2cdma_dat_entries_w\" -q sc2cdma_dat_entries");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2cdma_dat_updt <= 1'b0;
   end else begin
       sc2cdma_dat_updt <= dat_rls;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2cdma_dat_slices <= {14{1'b0}};
   end else begin
       if ((dat_rls) == 1'b1) begin
           sc2cdma_dat_slices <= sc2cdma_dat_slices_w[13:0];
       // VCS coverage off
       end else if ((dat_rls) == 1'b0) begin
       end else begin
           sc2cdma_dat_slices <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2cdma_dat_entries <= {15{1'b0}};
   end else begin
       if ((dat_rls) == 1'b1) begin
           sc2cdma_dat_entries <= sc2cdma_dat_entries_w;
       // VCS coverage off
       end else if ((dat_rls) == 1'b0) begin
       end else begin
           sc2cdma_dat_entries <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// input sg2dl package                                 /////
//////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////
///// generate data read sequence                        /////
//////////////////////////////////////////////////////////////
//: my $total_depth = 0 + 5;
//: my $wg_depth = 0;
//:
//: print "assign dl_in_pvld_d0 = sg2dl_pvld;\n";
//: print "assign dl_in_pd_d0 = sg2dl_pd;\n\n";
//:
//: for(my $i = 0; $i < $total_depth; $i ++) {
//: my $j = $i + 1;
//: &eperl::flop("-wid 1    -rval \"1'b0\"                                 -d \"dl_in_pvld_d${i}\" -q dl_in_pvld_d${j}");
//: &eperl::flop("-wid 31   -rval \"{31{1'b0}}\"  -en \"dl_in_pvld_d${i}\" -d \"dl_in_pd_d${i}\"   -q dl_in_pd_d${j}");
//: }
//:
//: my $d0 = $total_depth;
//: my $d1 = $wg_depth;
//:
//: print "assign dl_in_pvld = (is_winograd_d1[0]) ? dl_in_pvld_d${d1} : dl_in_pvld_d${d0};\n";
//: print "assign dl_in_pd = (is_winograd_d1[1]) ? dl_in_pd_d${d1} : dl_in_pd_d${d0};\n\n";
//: my $pipe_depth = 4;
//: my $i;
//: my $j;
//: print "assign dl_pvld_d0 = dl_in_pvld;\n";
//: print "assign dl_pd_d0 = dl_in_pd;\n\n";
//: for($i = 0; $i < $pipe_depth; $i ++) {
//: $j = $i + 1;
//: &eperl::flop("-nodeclare -rval \"1'b0\"                              -d \"dl_pvld_d${i}\"   -q dl_pvld_d${j}");
//: &eperl::flop("-nodeclare -rval \"{31{1'b0}}\"  -en \"dl_pvld_d${i}\" -d \"dl_pd_d${i}\"     -q dl_pd_d${j}");
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dl_in_pvld_d0 = sg2dl_pvld;
assign dl_in_pd_d0 = sg2dl_pd;

reg  dl_in_pvld_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d1 <= 1'b0;
   end else begin
       dl_in_pvld_d1 <= dl_in_pvld_d0;
   end
end
reg [30:0] dl_in_pd_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d1 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d0) == 1'b1) begin
           dl_in_pd_d1 <= dl_in_pd_d0;
       // VCS coverage off
       end else if ((dl_in_pvld_d0) == 1'b0) begin
       end else begin
           dl_in_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d2 <= 1'b0;
   end else begin
       dl_in_pvld_d2 <= dl_in_pvld_d1;
   end
end
reg [30:0] dl_in_pd_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d2 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d1) == 1'b1) begin
           dl_in_pd_d2 <= dl_in_pd_d1;
       // VCS coverage off
       end else if ((dl_in_pvld_d1) == 1'b0) begin
       end else begin
           dl_in_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d3 <= 1'b0;
   end else begin
       dl_in_pvld_d3 <= dl_in_pvld_d2;
   end
end
reg [30:0] dl_in_pd_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d3 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d2) == 1'b1) begin
           dl_in_pd_d3 <= dl_in_pd_d2;
       // VCS coverage off
       end else if ((dl_in_pvld_d2) == 1'b0) begin
       end else begin
           dl_in_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d4 <= 1'b0;
   end else begin
       dl_in_pvld_d4 <= dl_in_pvld_d3;
   end
end
reg [30:0] dl_in_pd_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d4 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d3) == 1'b1) begin
           dl_in_pd_d4 <= dl_in_pd_d3;
       // VCS coverage off
       end else if ((dl_in_pvld_d3) == 1'b0) begin
       end else begin
           dl_in_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dl_in_pvld_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pvld_d5 <= 1'b0;
   end else begin
       dl_in_pvld_d5 <= dl_in_pvld_d4;
   end
end
reg [30:0] dl_in_pd_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_in_pd_d5 <= {31{1'b0}};
   end else begin
       if ((dl_in_pvld_d4) == 1'b1) begin
           dl_in_pd_d5 <= dl_in_pd_d4;
       // VCS coverage off
       end else if ((dl_in_pvld_d4) == 1'b0) begin
       end else begin
           dl_in_pd_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
assign dl_in_pvld = (is_winograd_d1[0]) ? dl_in_pvld_d0 : dl_in_pvld_d5;
assign dl_in_pd = (is_winograd_d1[1]) ? dl_in_pd_d0 : dl_in_pd_d5;

assign dl_pvld_d0 = dl_in_pvld;
assign dl_pd_d0 = dl_in_pd;

always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d1 <= 1'b0;
   end else begin
       dl_pvld_d1 <= dl_pvld_d0;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d1 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d0) == 1'b1) begin
           dl_pd_d1 <= dl_pd_d0;
       // VCS coverage off
       end else if ((dl_pvld_d0) == 1'b0) begin
       end else begin
           dl_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d2 <= 1'b0;
   end else begin
       dl_pvld_d2 <= dl_pvld_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d2 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d1) == 1'b1) begin
           dl_pd_d2 <= dl_pd_d1;
       // VCS coverage off
       end else if ((dl_pvld_d1) == 1'b0) begin
       end else begin
           dl_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d3 <= 1'b0;
   end else begin
       dl_pvld_d3 <= dl_pvld_d2;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d3 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d2) == 1'b1) begin
           dl_pd_d3 <= dl_pd_d2;
       // VCS coverage off
       end else if ((dl_pvld_d2) == 1'b0) begin
       end else begin
           dl_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pvld_d4 <= 1'b0;
   end else begin
       dl_pvld_d4 <= dl_pvld_d3;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_pd_d4 <= {31{1'b0}};
   end else begin
       if ((dl_pvld_d3) == 1'b1) begin
           dl_pd_d4 <= dl_pd_d3;
       // VCS coverage off
       end else if ((dl_pvld_d3) == 1'b0) begin
       end else begin
           dl_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dl_pvld = (sub_h_total_g0[2] & dl_pvld_d1) |
                 (sub_h_total_g0[1] & dl_pvld_d3) |
                 (sub_h_total_g0[0] & dl_pvld_d4);
assign dl_pd = ({31 {sub_h_total_g1[2]}} & dl_pd_d1) |
               ({31 {sub_h_total_g1[1]}} & dl_pd_d3) |
               ({31 {sub_h_total_g1[0]}} & dl_pd_d4);
// PKT_UNPACK_WIRE( csc_dat_pkg , dl_ , dl_pd )
assign dl_w_offset[4:0] = dl_pd[4:0]; //this is weight offset
assign dl_h_offset[4:0] = dl_pd[9:5]; //weight offset
assign dl_channel_size[6:0] = dl_pd[16:10];
assign dl_stripe_length[6:0]= dl_pd[23:17];
assign dl_cur_sub_h[1:0] = dl_pd[25:24];
assign dl_block_end = dl_pd[26];
assign dl_channel_end = dl_pd[27];
assign dl_group_end = dl_pd[28];
assign dl_layer_end = dl_pd[29];
assign dl_dat_release = dl_pd[30];
////////////////////////// batch up counter //////////////////////////
assign {mon_batch_cnt_w,batch_cnt_w} = layer_st ? 6'b0 : is_batch_end ? 6'b0 : batch_cnt + 1'b1;
assign is_batch_end = (batch_cnt == batch_cmp);
//: &eperl::flop("-nodeclare   -rval \"{5{1'b0}}\"  -en \"layer_st | dat_exec_valid\" -d \"batch_cnt_w\" -q batch_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       batch_cnt <= {5{1'b0}};
   end else begin
       if ((layer_st | dat_exec_valid) == 1'b1) begin
           batch_cnt <= batch_cnt_w;
       // VCS coverage off
       end else if ((layer_st | dat_exec_valid) == 1'b0) begin
       end else begin
           batch_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// sub height up counter //////////////////////////
assign sub_h_cnt_inc = sub_h_cnt + 1'b1;
assign sub_h_cnt_w = (layer_st | is_sub_h_end) ? 2'b0 : sub_h_cnt_inc[1:0];
assign is_sub_h_end = (sub_h_cnt_inc == sub_h_cmp_g0);
assign sub_h_cnt_reg_en = layer_st | ((is_winograd_d1[2] | (|reg2dp_y_extension)) & dat_exec_valid);
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"sub_h_cnt_reg_en\" -d \"sub_h_cnt_w\" -q sub_h_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sub_h_cnt <= {2{1'b0}};
   end else begin
       if ((sub_h_cnt_reg_en) == 1'b1) begin
           sub_h_cnt <= sub_h_cnt_w;
       // VCS coverage off
       end else if ((sub_h_cnt_reg_en) == 1'b0) begin
       end else begin
           sub_h_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// stripe up counter //////////////////////////
assign {mon_stripe_cnt_inc,stripe_cnt_inc} = stripe_cnt + 1'b1;
assign stripe_cnt_w = layer_st ? 7'b0 :
                      (is_stripe_equal & ~is_sub_h_end) ? stripe_cnt :
                      is_stripe_end ? 7'b0 :
                      stripe_cnt_inc;
assign is_stripe_equal = is_batch_end & (stripe_cnt_inc == dl_stripe_length);
assign is_stripe_end = is_stripe_equal & is_sub_h_end;
assign stripe_cnt_reg_en = layer_st | (dat_exec_valid & is_batch_end);
//: &eperl::flop("-nodeclare   -rval \"{7{1'b0}}\"  -en \"stripe_cnt_reg_en\" -d \"stripe_cnt_w\" -q stripe_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       stripe_cnt <= {7{1'b0}};
   end else begin
       if ((stripe_cnt_reg_en) == 1'b1) begin
           stripe_cnt <= stripe_cnt_w;
       // VCS coverage off
       end else if ((stripe_cnt_reg_en) == 1'b0) begin
       end else begin
           stripe_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// pipe valid generator //////////////////////////
assign dat_pipe_local_valid_w = (dat_pipe_valid & is_stripe_equal) ? 1'b0 : dl_pvld ? 1'b1 : dat_pipe_local_valid;
assign dat_pipe_valid = dl_pvld | dat_pipe_local_valid;
assign dat_exec_valid = dl_pvld ? 1'b1 : (~(|stripe_cnt) & ~(|sub_h_cnt) & ~(|batch_cnt)) ? 1'b0 : dat_exec_valid_d1;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_pipe_local_valid_w\" -q dat_pipe_local_valid");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_pipe_valid\" -q dat_pipe_valid_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_exec_valid\" -q dat_exec_valid_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_pipe_local_valid <= 1'b0;
   end else begin
       dat_pipe_local_valid <= dat_pipe_local_valid_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_pipe_valid_d1 <= 1'b0;
   end else begin
       dat_pipe_valid_d1 <= dat_pipe_valid;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_exec_valid_d1 <= 1'b0;
   end else begin
       dat_exec_valid_d1 <= dat_exec_valid;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// request bytes //////////////////////////
assign dat_req_bytes = {1'b0, dl_channel_size};
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"dat_exec_valid\" -d \"dat_req_bytes\" -q dat_req_bytes_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_bytes_d1 <= {8{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_bytes_d1 <= dat_req_bytes;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_bytes_d1 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// output width coordinate counter //////////////////////////
// sub_h T, output will compute sub_h point in w direction
assign dataout_w_add = sub_h_cmp_g1;
assign {mon_dataout_w_cnt_inc,dataout_w_cnt_inc} = dataout_w_cnt + dataout_w_add;
assign is_w_end = is_batch_end & is_sub_h_end & (dataout_w_cnt >= dataout_width_cmp);
assign is_w_end_ahead = is_batch_end & (dataout_w_cnt >= dataout_width_cmp);
assign dataout_w_cnt_w = layer_st ? dataout_w_init :
                         (is_stripe_end & ~dl_channel_end) ? dataout_w_ori :
                         is_w_end ? dataout_w_init :
                         dataout_w_cnt_inc;
assign dataout_w_cnt_reg_en = layer_st | (dat_exec_valid & is_batch_end & is_sub_h_end);
assign dataout_w_ori_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_channel_end);
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"dataout_w_cnt_reg_en\" -d \"dataout_w_cnt_w\" -q dataout_w_cnt");
//: &eperl::flop("-nodeclare   -rval \"{13{1'b0}}\"  -en \"dataout_w_ori_reg_en\" -d \"dataout_w_cnt_w\" -q dataout_w_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dataout_w_cnt <= {13{1'b0}};
   end else begin
       if ((dataout_w_cnt_reg_en) == 1'b1) begin
           dataout_w_cnt <= dataout_w_cnt_w;
       // VCS coverage off
       end else if ((dataout_w_cnt_reg_en) == 1'b0) begin
       end else begin
           dataout_w_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dataout_w_ori <= {13{1'b0}};
   end else begin
       if ((dataout_w_ori_reg_en) == 1'b1) begin
           dataout_w_ori <= dataout_w_cnt_w;
       // VCS coverage off
       end else if ((dataout_w_ori_reg_en) == 1'b0) begin
       end else begin
           dataout_w_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// input channel coordinate counter, only feature  //////////////////////////
assign {mon_datain_c_cnt_inc,datain_c_cnt_inc} = datain_c_cnt + 1'b1;
assign is_last_channel = (datain_c_cnt == datain_channel_cmp);
assign datain_c_cnt_w = layer_st ? 11'b0 : dl_channel_end ? 11'b0 : datain_c_cnt_inc;
assign datain_c_cnt_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_block_end);
//: &eperl::flop("-nodeclare   -rval \"{11{1'b0}}\"  -en \"datain_c_cnt_reg_en\" -d \"datain_c_cnt_w\" -q datain_c_cnt");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_c_cnt <= {11{1'b0}};
   end else begin
       if ((datain_c_cnt_reg_en) == 1'b1) begin
           datain_c_cnt <= datain_c_cnt_w;
       // VCS coverage off
       end else if ((datain_c_cnt_reg_en) == 1'b0) begin
       end else begin
           datain_c_cnt <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// input width coordinate counter, feature/image dedicated counter //////////////////////////
assign datain_w_cnt_st = (is_img) ? 14'b0 : (is_winograd) ? 14'h2 : 13'b0 - reg2dp_pad_left;
assign {mon_datain_w_cnt_inc,datain_w_cnt_inc} = (is_winograd_d1[3]) ? (datain_w_cnt + 2'h2) : (datain_w_cnt + conv_x_stride);
//full data cube w counter,start form negtive, only for feature data. non-image, by element
assign datain_w_cnt_w = layer_st ? datain_w_cnt_st :
                        (is_stripe_end & ~dl_channel_end) ? datain_w_ori :
                        is_w_end ? datain_w_cnt_st :
                        datain_w_cnt_inc;
assign dl_w_offset_ext = dl_w_offset * x_dilate;
assign {mon_datain_w_cur,datain_w_cur} = datain_w_cnt + dl_w_offset_ext; //by element
assign datain_w_cnt_reg_en = layer_st | (dat_exec_valid & is_batch_end & is_sub_h_end & ~is_img_d1[0]);
assign datain_w_ori_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_channel_end & ~is_img_d1[1]);
//notice:after sub_h T, pixel_x_add elements in W direction is used by CMAC
assign pixel_x_cnt_add = (is_sub_h_end) ? pixel_x_add : 6'b0;
//assign {mon_pixel_w_cnt_w,pixel_w_cnt_w} = (layer_st_d1) ? {{11{1'b0}}, pixel_x_init} :
// (is_stripe_end & dl_block_end & dl_channel_end & is_w_end) ? {{11{1'b0}}, pixel_x_init} :
// (is_stripe_end & dl_block_end & dl_channel_end & ~is_w_end) ? (pixel_w_ch_ori + pixel_ch_stride) :
// (is_stripe_end & dl_block_end & ~dl_channel_end) ? (pixel_w_ch_ori + pixel_x_init_offset) :
// (is_stripe_end & ~dl_block_end) ? {1'b0, pixel_w_ori} :
// (pixel_w_cnt + pixel_x_cnt_add);
//channel count.
wire [12:0] total_channel_op = (reg2dp_weight_channel_ext[6 -1:0]=={6{1'b0}}) ?
                        reg2dp_weight_channel_ext[12:6] : reg2dp_weight_channel_ext[12:6]+1'b1;
reg [12:0] channel_op_cnt;
wire mon_channel_op_cnt_nxt;
wire [12:0] channel_op_cnt_nxt;
assign {mon_channel_op_cnt_nxt, channel_op_cnt_nxt} = dl_channel_end&is_stripe_end ? 13'h2 :
                                                        dl_block_end&is_stripe_end ? channel_op_cnt + 1'b1 :
                                                        channel_op_cnt;
//: &eperl::flop("-q channel_op_cnt  -d \"channel_op_cnt_nxt\"  -wid 13  -rval \"13'h2\" -nodeclare ");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       channel_op_cnt <= 13'h2;
   end else begin
       channel_op_cnt <= channel_op_cnt_nxt;
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
wire next_is_last_channel = (channel_op_cnt >= total_channel_op);
//notice, after pre-extention, image weight w_total <=128
assign {mon_pixel_w_cnt_w,pixel_w_cnt_w} = (layer_st_d1) ? {{11{1'b0}}, pixel_x_init} :
                        (is_stripe_end & dl_block_end & dl_channel_end & is_w_end) ? {{11{1'b0}}, pixel_x_init} :
                        (is_stripe_end & dl_block_end & dl_channel_end & ~is_w_end) ? (pixel_w_ch_ori + pixel_ch_stride) :
//(is_stripe_end & dl_block_end & ~dl_channel_end) ? (pixel_w_ori + dl_in_pd_d0[16:10]) :
                        (is_stripe_end & dl_block_end & next_is_last_channel) ? (pixel_w_ori + pixel_x_init_offset) :
                        (is_stripe_end & dl_block_end & ~next_is_last_channel) ? (pixel_w_ori + 8'h40  ) :
                        (is_stripe_end & ~dl_block_end) ? {1'b0, pixel_w_ori} :
                        (pixel_w_cnt + pixel_x_cnt_add);
assign pixel_w_cur = {{6 -1{1'b0}},pixel_w_cnt[15:6]}; //by entry 
assign pixel_w_cnt_reg_en = layer_st_d1 | (dat_exec_valid & is_img_d1[2] & (is_sub_h_end | is_w_end));
assign pixel_w_ori_reg_en = layer_st_d1 | (dat_exec_valid & is_img_d1[3] & is_stripe_end & dl_block_end);
assign pixel_ch_ori_reg_en = layer_st_d1 | (dat_exec_valid & is_img_d1[4] & is_stripe_end & dl_block_end & dl_channel_end);
assign pixel_force_fetch = (is_img_d1[0] & dat_req_stripe_st) ? 1'b1 : (pixel_force_clr_d1) ? 1'b0 : pixel_force_fetch_d1;
assign pixel_force_clr = is_img_d1[0] & is_sub_h_end & (pixel_force_fetch | pixel_force_fetch_d1);
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_w_cnt_reg_en\" -d \"datain_w_cnt_w\" -q datain_w_cnt");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_w_ori_reg_en\" -d \"datain_w_cnt_w\" -q datain_w_ori");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"pixel_w_cnt_reg_en\" -d \"pixel_w_cnt_w\" -q pixel_w_cnt");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"pixel_w_ori_reg_en\" -d \"pixel_w_cnt_w\" -q pixel_w_ori");
//: &eperl::flop("-nodeclare   -rval \"{16{1'b0}}\"  -en \"pixel_ch_ori_reg_en\" -d \"pixel_w_cnt_w\" -q pixel_w_ch_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_w_cnt <= {14{1'b0}};
   end else begin
       if ((datain_w_cnt_reg_en) == 1'b1) begin
           datain_w_cnt <= datain_w_cnt_w;
       // VCS coverage off
       end else if ((datain_w_cnt_reg_en) == 1'b0) begin
       end else begin
           datain_w_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_w_ori <= {14{1'b0}};
   end else begin
       if ((datain_w_ori_reg_en) == 1'b1) begin
           datain_w_ori <= datain_w_cnt_w;
       // VCS coverage off
       end else if ((datain_w_ori_reg_en) == 1'b0) begin
       end else begin
           datain_w_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_w_cnt <= {16{1'b0}};
   end else begin
       if ((pixel_w_cnt_reg_en) == 1'b1) begin
           pixel_w_cnt <= pixel_w_cnt_w;
       // VCS coverage off
       end else if ((pixel_w_cnt_reg_en) == 1'b0) begin
       end else begin
           pixel_w_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_w_ori <= {16{1'b0}};
   end else begin
       if ((pixel_w_ori_reg_en) == 1'b1) begin
           pixel_w_ori <= pixel_w_cnt_w;
       // VCS coverage off
       end else if ((pixel_w_ori_reg_en) == 1'b0) begin
       end else begin
           pixel_w_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_w_ch_ori <= {16{1'b0}};
   end else begin
       if ((pixel_ch_ori_reg_en) == 1'b1) begin
           pixel_w_ch_ori <= pixel_w_cnt_w;
       // VCS coverage off
       end else if ((pixel_ch_ori_reg_en) == 1'b0) begin
       end else begin
           pixel_w_ch_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// input height coordinate counter, feature/image both  //////////////////////////
// full data cube h counter, start form negative
assign datain_h_cnt_st = (is_winograd) ? 14'b0 : 14'b0 - reg2dp_pad_top;
assign {mon_datain_h_cnt_inc, datain_h_cnt_inc} = datain_h_cnt + conv_y_stride;
assign datain_h_cnt_w = (layer_st | (is_stripe_end & dl_group_end)) ? datain_h_cnt_st :
                        (is_stripe_end & ~dl_channel_end) ? datain_h_ori :
                        is_w_end ? datain_h_cnt_inc :
                        datain_h_cnt;
assign datain_h_cnt_reg_en = layer_st | (dat_exec_valid & ((is_stripe_end & ~dl_channel_end) | is_w_end));
assign datain_h_ori_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_channel_end);
assign dl_h_offset_ext = dl_h_offset * y_dilate;
assign {mon_datain_h_cur,datain_h_cur} = datain_h_cnt + dl_h_offset_ext + sub_h_cnt;
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_h_cnt_reg_en\" -d \"datain_h_cnt_w\" -q datain_h_cnt");
//: &eperl::flop("-nodeclare   -rval \"{14{1'b0}}\"  -en \"datain_h_ori_reg_en\" -d \"datain_h_cnt_w\" -q datain_h_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_h_cnt <= {14{1'b0}};
   end else begin
       if ((datain_h_cnt_reg_en) == 1'b1) begin
           datain_h_cnt <= datain_h_cnt_w;
       // VCS coverage off
       end else if ((datain_h_cnt_reg_en) == 1'b0) begin
       end else begin
           datain_h_cnt <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       datain_h_ori <= {14{1'b0}};
   end else begin
       if ((datain_h_ori_reg_en) == 1'b1) begin
           datain_h_ori <= datain_h_cnt_w;
       // VCS coverage off
       end else if ((datain_h_ori_reg_en) == 1'b0) begin
       end else begin
           datain_h_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// fetch valid generate //////////////////////////
assign dat_conv_req_dummy = (datain_w_cur[13 ]) | (datain_w_cur > {1'b0, datain_width_cmp})
                            | (datain_h_cur[13 ]) | (datain_h_cur > {1'b0, datain_height_cmp});
assign dat_wg_req_dummy = 1'b0;
assign dat_wg_req_skip = ((|datain_w_cur[13:2]) & datain_w_cur[1] & (|stripe_cnt[6:1]));
assign dat_img_req_dummy = (datain_h_cur[13]) | (datain_h_cur > {1'b0, datain_height_cmp});
//w address(in entry) is bigger than avilable entrys
assign dat_img_req_skip = ({{15 -12{1'b0}},w_bias_w[13:2]} > entries_cmp[15 -1:0]);
assign dat_req_dummy = is_img_d1[5] ? dat_img_req_dummy : is_winograd_d1[4] ? dat_wg_req_dummy : dat_conv_req_dummy;
assign dat_req_skip = (is_winograd_d1[5] & dat_wg_req_skip) | (is_img_d1[6] & dat_img_req_skip);
assign dat_req_valid = (dat_exec_valid & ~dat_req_dummy & ~dat_req_skip);
//Add corner case
assign dat_req_sub_c_w = ~is_img_d1[7] ? datain_c_cnt[0] : dl_block_end;
assign dat_req_sub_w_w = is_winograd_d1[6] ? {1'b0, ~datain_w_cur[1]} : datain_w_cur[1:0];
assign dat_req_sub_w_st_en = dat_exec_valid & (sub_h_cnt == 2'h0);
assign dat_req_batch_index = batch_cnt;
assign dat_req_stripe_st = dl_pvld;
assign dat_req_stripe_end = is_stripe_equal & dat_pipe_valid;
assign dat_req_channel_end = dl_channel_end;
assign dat_req_layer_end = dl_layer_end;
// PKT_PACK_WIRE( nvdla_stripe_info , dat_req_ , dat_req_flag_w )
assign dat_req_flag_w[4:0] = dat_req_batch_index[4:0];
assign dat_req_flag_w[5] = dat_req_stripe_st ;
assign dat_req_flag_w[6] = dat_req_stripe_end ;
assign dat_req_flag_w[7] = dat_req_channel_end ;
assign dat_req_flag_w[8] = dat_req_layer_end ;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_req_valid\" -q dat_req_valid_d1");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid\" -d \"dat_req_sub_w_w\" -q dat_req_sub_w_d1");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid\" -d \"sub_h_cnt\" -q dat_req_sub_h_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"dat_req_sub_c_w\" -q dat_req_sub_c_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"is_last_channel\" -q dat_req_ch_end_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"dat_req_dummy\" -q dat_req_dummy_d1");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid\" -d \"dl_cur_sub_h\" -q dat_req_cur_sub_h_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_req_sub_w_st_en\" -d \"dat_req_stripe_st\" -q dat_req_sub_w_st_d1");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_exec_valid\" -d \"dat_req_flag_w\" -q dat_req_flag_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"dl_dat_release & is_stripe_equal & dat_pipe_valid\" -q dat_req_rls_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"pixel_force_fetch\" -q pixel_force_fetch_d1");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid\" -d \"pixel_force_clr\" -q pixel_force_clr_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_valid_d1 <= 1'b0;
   end else begin
       dat_req_valid_d1 <= dat_req_valid;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_d1 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_sub_w_d1 <= dat_req_sub_w_w;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_sub_w_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_d1 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_sub_h_d1 <= sub_h_cnt;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_sub_h_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_c_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_sub_c_d1 <= dat_req_sub_c_w;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_sub_c_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_ch_end_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_ch_end_d1 <= is_last_channel;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_ch_end_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_dummy_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_dummy_d1 <= dat_req_dummy;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_dummy_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_cur_sub_h_d1 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_cur_sub_h_d1 <= dl_cur_sub_h;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_cur_sub_h_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_st_d1 <= 1'b0;
   end else begin
       if ((dat_req_sub_w_st_en) == 1'b1) begin
           dat_req_sub_w_st_d1 <= dat_req_stripe_st;
       // VCS coverage off
       end else if ((dat_req_sub_w_st_en) == 1'b0) begin
       end else begin
           dat_req_sub_w_st_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_flag_d1 <= {9{1'b0}};
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_flag_d1 <= dat_req_flag_w;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_flag_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_rls_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           dat_req_rls_d1 <= dl_dat_release & is_stripe_equal & dat_pipe_valid;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           dat_req_rls_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_force_fetch_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           pixel_force_fetch_d1 <= pixel_force_fetch;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           pixel_force_fetch_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       pixel_force_clr_d1 <= 1'b0;
   end else begin
       if ((dat_exec_valid) == 1'b1) begin
           pixel_force_clr_d1 <= pixel_force_clr;
       // VCS coverage off
       end else if ((dat_exec_valid) == 1'b0) begin
       end else begin
           pixel_force_clr_d1 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// generate data read address                         /////
//////////////////////////////////////////////////////////////
////////////////////////// data read index generator: 1st stage //////////////////////////
//channel bias, by w_in element
//assign c_bias_add = (~is_img_d1[8] & datain_c_cnt[0]) ? datain_width[12 -1:0] : 12'b0;
assign c_bias_add = (~is_img_d1[8]) ? datain_width[12 -1:0] : 12'b0;
assign {mon_c_bias_w, c_bias_w} = layer_st ? 13'b0 : (is_stripe_end & dl_channel_end) ? 13'b0 : c_bias + c_bias_add;
assign c_bias_reg_en = layer_st | (dat_exec_valid & is_stripe_end & dl_block_end);
assign c_bias_d1_reg_en = (c_bias != c_bias_d1);
//height bias, by element
assign {mon_h_bias_0_w,h_bias_0_w} = datain_h_cnt[13:0] * h_bias_0_stride;
assign {mon_h_bias_1_w,h_bias_1_w} = dl_h_offset * h_bias_1_stride;
assign {mon_h_bias_2_w,h_bias_2_w} = batch_cnt * h_bias_2_stride;
assign {mon_h_bias_3_w,h_bias_3_w} = layer_st ? 13'b0 :sub_h_cnt * h_bias_3_stride;
assign h_bias_reg_en[0] = dat_exec_valid;
assign h_bias_reg_en[1] = layer_st | (dat_exec_valid & (is_winograd_d1[7] | is_img_d1[9]));
//width bias, by entry in image, by element in feature data

assign w_bias_int8 = is_img_d1[10] ? {pixel_w_cur} : //by entry in image 
                     is_winograd_d1[8] ? {1'b0, datain_w_cnt} :
                     (~is_last_channel | is_winograd_d1[8]) ? {2'b0,datain_w_cur[12:0]} ://not last channel, by element
                     (dat_req_bytes > 8'h20) ? {2'b0,datain_w_cur[12:0]} : //last channel & request >1/2*entry
                     {3'b0, datain_w_cur[12:1]}; //last channel & request<=1/2*entry

assign w_bias_int8 = is_img_d1[10] ? {pixel_w_cur} : //by entry in image 
                     is_winograd_d1[8] ? {1'b0, datain_w_cnt} :
                     (~is_last_channel | is_winograd_d1[8]) ? {2'b0,datain_w_cur[12:0]} ://not last channel, by element
                     (dat_req_bytes > 8'h20) ? {2'b0,datain_w_cur[12:0]} : //last channel & request >1/2*entry
                     (dat_req_bytes <= 8'h10) ? {4'b0, datain_w_cur[12:2]} : //last channel & request <=1/4*entry
                     {3'b0, datain_w_cur[12:1]}; //last channel & (1/4*entry<request<=1/2*entry)
assign w_bias_w = w_bias_int8[13:0];
assign w_bias_reg_en = dat_exec_valid;
assign dat_req_base_d1 = dat_entry_st[13 -1:0];
//: my $kk=13;
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"c_bias_reg_en\" -d \"c_bias_w\" -q c_bias");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"c_bias_d1_reg_en\" -d \"c_bias\" -q c_bias_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[0]\" -d \"h_bias_0_w\" -q h_bias_0_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[0]\" -d \"h_bias_1_w\" -q h_bias_1_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[0]\" -d \"h_bias_2_w\" -q h_bias_2_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"h_bias_reg_en[1]\" -d \"h_bias_3_w\" -q h_bias_3_d1");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"w_bias_reg_en\" -d \"w_bias_w\" -q w_bias_d1");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       c_bias <= {13{1'b0}};
   end else begin
       if ((c_bias_reg_en) == 1'b1) begin
           c_bias <= c_bias_w;
       // VCS coverage off
       end else if ((c_bias_reg_en) == 1'b0) begin
       end else begin
           c_bias <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       c_bias_d1 <= {13{1'b0}};
   end else begin
       if ((c_bias_d1_reg_en) == 1'b1) begin
           c_bias_d1 <= c_bias;
       // VCS coverage off
       end else if ((c_bias_d1_reg_en) == 1'b0) begin
       end else begin
           c_bias_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_0_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[0]) == 1'b1) begin
           h_bias_0_d1 <= h_bias_0_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[0]) == 1'b0) begin
       end else begin
           h_bias_0_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_1_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[0]) == 1'b1) begin
           h_bias_1_d1 <= h_bias_1_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[0]) == 1'b0) begin
       end else begin
           h_bias_1_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_2_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[0]) == 1'b1) begin
           h_bias_2_d1 <= h_bias_2_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[0]) == 1'b0) begin
       end else begin
           h_bias_2_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       h_bias_3_d1 <= {13{1'b0}};
   end else begin
       if ((h_bias_reg_en[1]) == 1'b1) begin
           h_bias_3_d1 <= h_bias_3_w;
       // VCS coverage off
       end else if ((h_bias_reg_en[1]) == 1'b0) begin
       end else begin
           h_bias_3_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       w_bias_d1 <= {13{1'b0}};
   end else begin
       if ((w_bias_reg_en) == 1'b1) begin
           w_bias_d1 <= w_bias_w;
       // VCS coverage off
       end else if ((w_bias_reg_en) == 1'b0) begin
       end else begin
           w_bias_d1 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
////////////////////////// data read index generator: 2st stage //////////////////////////
wire [13 -1:0] dat_req_addr_minus1;
wire mon_dat_req_addr_minus1;
wire is_dat_req_addr_minus1_wrap;
wire [13 -1:0] dat_req_addr_minus1_wrap;
wire [13 -1:0] dat_req_addr_minus1_real;
assign {mon_h_bias_d1,h_bias_d1} = h_bias_0_d1 + h_bias_1_d1 + h_bias_2_d1 + h_bias_3_d1;
//assign {mon_dat_req_addr_sum,dat_req_addr_sum} = dat_req_base_d1 + c_bias_d1 + h_bias_d1 + w_bias_d1; //by entry
assign dat_req_addr_sum = dat_req_base_d1 + c_bias_d1 + h_bias_d1 + w_bias_d1; //by entry
assign is_dat_req_addr_wrap = (dat_req_addr_sum >= {1'b0,data_bank, {9{1'b0}}});
assign {mon_dat_req_addr_wrap,dat_req_addr_wrap} = dat_req_addr_sum[13:0] - {1'b0,data_bank, {9{1'b0}}};
assign dat_req_addr_w = (layer_st | dat_req_dummy_d1) ? {13{1'b1}} : is_dat_req_addr_wrap ? dat_req_addr_wrap : dat_req_addr_sum[13 -1:0]; //get the adress sends to cbuf
assign {mon_dat_req_addr_minus1,dat_req_addr_minus1} = dat_req_addr_w-1'b1;
assign is_dat_req_addr_minus1_wrap = (dat_req_addr_minus1 >= {data_bank, {9{1'b0}}}); //only one case: 0-1=ffff would introduce wrap  
assign dat_req_addr_minus1_wrap = {data_bank, {9{1'b1}}};
assign dat_req_addr_minus1_real = is_dat_req_addr_minus1_wrap ? dat_req_addr_minus1_wrap : dat_req_addr_minus1;
assign sc2buf_dat_rd_en_w = dat_req_valid_d1 & ((dat_req_addr_last != dat_req_addr_w) | pixel_force_fetch_d1);
assign dat_req_addr_last = (dat_req_sub_h_d1 == 2'h0) ? dat_req_sub_h_0_addr :
                           (dat_req_sub_h_d1 == 2'h1) ? dat_req_sub_h_1_addr :
                           (dat_req_sub_h_d1 == 2'h2) ? dat_req_sub_h_2_addr :
                           dat_req_sub_h_3_addr;
assign dat_req_sub_h_0_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h0));
assign dat_req_sub_h_1_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h1));
assign dat_req_sub_h_2_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h2));
assign dat_req_sub_h_3_addr_en = layer_st | ((dat_req_valid_d1 | dat_req_dummy_d1) & (dat_req_sub_h_d1 == 2'h3));

wire [13 -1:0] sc2buf_dat_rd_addr_w;
assign sc2buf_dat_rd_addr_w = dat_req_addr_w;
//: my $kk=13;
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_0_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_0_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_1_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_1_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_2_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_2_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"dat_req_sub_h_3_addr_en\" -d \"dat_req_addr_w\" -q dat_req_sub_h_3_addr");
//: my $kk=13;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"sc2buf_dat_rd_en_w\" -q sc2buf_dat_rd_en");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"layer_st | sc2buf_dat_rd_en_w\" -d \"sc2buf_dat_rd_addr_w\" -q sc2buf_dat_rd_addr");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b1}}\"  -en \"layer_st | sc2buf_dat_rd_en_w\" -d \"sc2buf_dat_rd_next1_addr_w\" -q sc2buf_dat_rd_next1_addr");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_pipe_valid_d1\" -q dat_pipe_valid_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_exec_valid_d1\" -q dat_exec_valid_d2");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_w_d1\" -q dat_req_sub_w_d2");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_h_d1\" -q dat_req_sub_h_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_c_d1\" -q dat_req_sub_c_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_ch_end_d1\" -q dat_req_ch_end_d2");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_bytes_d1\" -q dat_req_bytes_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_dummy_d1\" -q dat_req_dummy_d2");
//: &eperl::flop("-nodeclare   -rval \"{2{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_cur_sub_h_d1\" -q dat_req_cur_sub_h_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_sub_w_st_d1\" -q dat_req_sub_w_st_d2");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"  -en \"dat_exec_valid_d1\" -d \"dat_req_rls_d1\" -q dat_req_rls_d2");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_exec_valid_d1\" -d \"dat_req_flag_d1\" -q dat_req_flag_d2");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_0_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_0_addr_en) == 1'b1) begin
           dat_req_sub_h_0_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_0_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_0_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_1_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_1_addr_en) == 1'b1) begin
           dat_req_sub_h_1_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_1_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_1_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_2_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_2_addr_en) == 1'b1) begin
           dat_req_sub_h_2_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_2_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_2_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_3_addr <= {13{1'b1}};
   end else begin
       if ((dat_req_sub_h_3_addr_en) == 1'b1) begin
           dat_req_sub_h_3_addr <= dat_req_addr_w;
       // VCS coverage off
       end else if ((dat_req_sub_h_3_addr_en) == 1'b0) begin
       end else begin
           dat_req_sub_h_3_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2buf_dat_rd_en <= 1'b0;
   end else begin
       sc2buf_dat_rd_en <= sc2buf_dat_rd_en_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2buf_dat_rd_addr <= {13{1'b1}};
   end else begin
       if ((layer_st | sc2buf_dat_rd_en_w) == 1'b1) begin
           sc2buf_dat_rd_addr <= sc2buf_dat_rd_addr_w;
       // VCS coverage off
       end else if ((layer_st | sc2buf_dat_rd_en_w) == 1'b0) begin
       end else begin
           sc2buf_dat_rd_addr <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_pipe_valid_d2 <= 1'b0;
   end else begin
       dat_pipe_valid_d2 <= dat_pipe_valid_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_exec_valid_d2 <= 1'b0;
   end else begin
       dat_exec_valid_d2 <= dat_exec_valid_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_d2 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_w_d2 <= dat_req_sub_w_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_w_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_h_d2 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_h_d2 <= dat_req_sub_h_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_h_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_c_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_c_d2 <= dat_req_sub_c_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_c_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_ch_end_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_ch_end_d2 <= dat_req_ch_end_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_ch_end_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_bytes_d2 <= {8{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_bytes_d2 <= dat_req_bytes_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_bytes_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_dummy_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_dummy_d2 <= dat_req_dummy_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_dummy_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_cur_sub_h_d2 <= {2{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_cur_sub_h_d2 <= dat_req_cur_sub_h_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_cur_sub_h_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_sub_w_st_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_sub_w_st_d2 <= dat_req_sub_w_st_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_sub_w_st_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_rls_d2 <= 1'b0;
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_rls_d2 <= dat_req_rls_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_rls_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_req_flag_d2 <= {9{1'b0}};
   end else begin
       if ((dat_exec_valid_d1) == 1'b1) begin
           dat_req_flag_d2 <= dat_req_flag_d1;
       // VCS coverage off
       end else if ((dat_exec_valid_d1) == 1'b0) begin
       end else begin
           dat_req_flag_d2 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// sideband pipeline                                  /////
//////////////////////////////////////////////////////////////
assign dat_req_pipe_pvld = dat_pipe_valid_d2;
assign dat_req_pipe_sub_w = dat_req_sub_w_d2;
assign dat_req_pipe_sub_h = dat_req_sub_h_d2;
assign dat_req_pipe_sub_c = dat_req_sub_c_d2;
assign dat_req_pipe_ch_end = dat_req_ch_end_d2;
assign dat_req_pipe_bytes = dat_req_bytes_d2;
assign dat_req_pipe_dummy = dat_req_dummy_d2;
assign dat_req_pipe_cur_sub_h = dat_req_cur_sub_h_d2;
assign dat_req_pipe_sub_w_st = dat_req_sub_w_st_d2;
assign dat_req_pipe_rls = dat_req_rls_d2;
assign dat_req_pipe_flag = dat_req_flag_d2;
assign dat_req_exec_pvld = dat_exec_valid_d2;
assign dat_req_exec_dummy = dat_req_dummy_d2;
assign dat_req_exec_sub_h = dat_req_sub_h_d2;
// PKT_PACK_WIRE( csc_dat_req_pkg , dat_req_pipe_ , dat_req_pipe_pd )
assign dat_req_pipe_pd[1:0] = dat_req_pipe_sub_w[1:0];
assign dat_req_pipe_pd[3:2] = dat_req_pipe_sub_h[1:0];
assign dat_req_pipe_pd[4] = dat_req_pipe_sub_c ;
assign dat_req_pipe_pd[5] = dat_req_pipe_ch_end ;
assign dat_req_pipe_pd[6] = 1'b0 ;
assign dat_req_pipe_pd[14:7] = dat_req_pipe_bytes[7:0];
assign dat_req_pipe_pd[16:15] = dat_req_pipe_cur_sub_h[1:0];
assign dat_req_pipe_pd[17] = dat_req_pipe_dummy ;
assign dat_req_pipe_pd[18] = dat_req_pipe_sub_w_st ;
assign dat_req_pipe_pd[19] = dat_req_pipe_rls ;
assign dat_req_pipe_pd[28:20] = dat_req_pipe_flag[8:0];
//add latency for data request contorl signal
//: my $pipe_depth = 6;
//: my $i;
//: my $j;
//: if($pipe_depth == 0) {
//: print "assign dat_rsp_pipe_pvld = dat_req_pipe_pvld;\n";
//: print "assign dat_rsp_pipe_pd = dat_req_pipe_pd;\n";
//: print "assign dat_rsp_exec_pvld = dat_req_exec_pvld;\n";
//: print "assign dat_rsp_exec_dummy = dat_req_exec_dummy;\n";
//: print "assign dat_rsp_exec_sub_h = dat_req_exec_sub_h;\n\n";
//: } else {
//: print "assign dat_rsp_pipe_pvld_d0 = dat_req_pipe_pvld;\n";
//: print "assign dat_rsp_pipe_pd_d0 = dat_req_pipe_pd;\n";
//: print "assign dat_rsp_exec_pvld_d0 = dat_req_exec_pvld;\n";
//: print "assign dat_rsp_exec_dummy_d0 = dat_req_exec_dummy;\n";
//: print "assign dat_rsp_exec_sub_h_d0 = dat_req_exec_sub_h;\n\n";
//: for($i = 0; $i < $pipe_depth; $i ++) {
//: $j = $i + 1;
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -d \"dat_rsp_pipe_pvld_d${i}\"  -q dat_rsp_pipe_pvld_d${j}");
//: &eperl::flop("-wid 29  -rval \"{29{1'b0}}\" -en \"dat_rsp_pipe_pvld_d${i}\" -d \"dat_rsp_pipe_pd_d${i}\"    -q dat_rsp_pipe_pd_d${j}");
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -d \"dat_rsp_exec_pvld_d${i}\"  -q dat_rsp_exec_pvld_d${j}");
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -en \"dat_rsp_exec_pvld_d${i}\" -d \"dat_rsp_exec_dummy_d${i}\" -q dat_rsp_exec_dummy_d${j}");
//: &eperl::flop("-wid 2   -rval \"{2{1'b0}}\"  -en \"dat_rsp_exec_pvld_d${i}\" -d \"dat_rsp_exec_sub_h_d${i}\" -q dat_rsp_exec_sub_h_d${j}");
//: }
//: print "assign dat_rsp_pipe_pvld = dat_rsp_pipe_pvld_d${i};\n";
//: print "assign dat_rsp_pipe_pd = dat_rsp_pipe_pd_d${i};\n";
//: print "assign dat_rsp_exec_pvld = dat_rsp_exec_pvld_d${i};\n";
//: print "assign dat_rsp_exec_dummy = dat_rsp_exec_dummy_d${i};\n";
//: print "assign dat_rsp_exec_sub_h = dat_rsp_exec_sub_h_d${i};\n\n";
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_rsp_pipe_pvld_d0 = dat_req_pipe_pvld;
assign dat_rsp_pipe_pd_d0 = dat_req_pipe_pd;
assign dat_rsp_exec_pvld_d0 = dat_req_exec_pvld;
assign dat_rsp_exec_dummy_d0 = dat_req_exec_dummy;
assign dat_rsp_exec_sub_h_d0 = dat_req_exec_sub_h;

reg  dat_rsp_pipe_pvld_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d1 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d1 <= dat_rsp_pipe_pvld_d0;
   end
end
reg [28:0] dat_rsp_pipe_pd_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d1 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d0) == 1'b1) begin
           dat_rsp_pipe_pd_d1 <= dat_rsp_pipe_pd_d0;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d1 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d1 <= dat_rsp_exec_pvld_d0;
   end
end
reg  dat_rsp_exec_dummy_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d1 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d0) == 1'b1) begin
           dat_rsp_exec_dummy_d1 <= dat_rsp_exec_dummy_d0;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d1 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d0) == 1'b1) begin
           dat_rsp_exec_sub_h_d1 <= dat_rsp_exec_sub_h_d0;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d2 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d2 <= dat_rsp_pipe_pvld_d1;
   end
end
reg [28:0] dat_rsp_pipe_pd_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d2 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d1) == 1'b1) begin
           dat_rsp_pipe_pd_d2 <= dat_rsp_pipe_pd_d1;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d2 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d2 <= dat_rsp_exec_pvld_d1;
   end
end
reg  dat_rsp_exec_dummy_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d2 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d1) == 1'b1) begin
           dat_rsp_exec_dummy_d2 <= dat_rsp_exec_dummy_d1;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d2 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d1) == 1'b1) begin
           dat_rsp_exec_sub_h_d2 <= dat_rsp_exec_sub_h_d1;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d3 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d3 <= dat_rsp_pipe_pvld_d2;
   end
end
reg [28:0] dat_rsp_pipe_pd_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d3 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d2) == 1'b1) begin
           dat_rsp_pipe_pd_d3 <= dat_rsp_pipe_pd_d2;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d3 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d3 <= dat_rsp_exec_pvld_d2;
   end
end
reg  dat_rsp_exec_dummy_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d3 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d2) == 1'b1) begin
           dat_rsp_exec_dummy_d3 <= dat_rsp_exec_dummy_d2;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d3 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d2) == 1'b1) begin
           dat_rsp_exec_sub_h_d3 <= dat_rsp_exec_sub_h_d2;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d4 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d4 <= dat_rsp_pipe_pvld_d3;
   end
end
reg [28:0] dat_rsp_pipe_pd_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d4 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d3) == 1'b1) begin
           dat_rsp_pipe_pd_d4 <= dat_rsp_pipe_pd_d3;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d4 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d4 <= dat_rsp_exec_pvld_d3;
   end
end
reg  dat_rsp_exec_dummy_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d4 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d3) == 1'b1) begin
           dat_rsp_exec_dummy_d4 <= dat_rsp_exec_dummy_d3;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d4 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d3) == 1'b1) begin
           dat_rsp_exec_sub_h_d4 <= dat_rsp_exec_sub_h_d3;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d5 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d5 <= dat_rsp_pipe_pvld_d4;
   end
end
reg [28:0] dat_rsp_pipe_pd_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d5 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d4) == 1'b1) begin
           dat_rsp_pipe_pd_d5 <= dat_rsp_pipe_pd_d4;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d4) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d5 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d5 <= dat_rsp_exec_pvld_d4;
   end
end
reg  dat_rsp_exec_dummy_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d5 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d4) == 1'b1) begin
           dat_rsp_exec_dummy_d5 <= dat_rsp_exec_dummy_d4;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d4) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d5 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d4) == 1'b1) begin
           dat_rsp_exec_sub_h_d5 <= dat_rsp_exec_sub_h_d4;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d4) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d5 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_pipe_pvld_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pvld_d6 <= 1'b0;
   end else begin
       dat_rsp_pipe_pvld_d6 <= dat_rsp_pipe_pvld_d5;
   end
end
reg [28:0] dat_rsp_pipe_pd_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pipe_pd_d6 <= {29{1'b0}};
   end else begin
       if ((dat_rsp_pipe_pvld_d5) == 1'b1) begin
           dat_rsp_pipe_pd_d6 <= dat_rsp_pipe_pd_d5;
       // VCS coverage off
       end else if ((dat_rsp_pipe_pvld_d5) == 1'b0) begin
       end else begin
           dat_rsp_pipe_pd_d6 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_rsp_exec_pvld_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_pvld_d6 <= 1'b0;
   end else begin
       dat_rsp_exec_pvld_d6 <= dat_rsp_exec_pvld_d5;
   end
end
reg  dat_rsp_exec_dummy_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_dummy_d6 <= 1'b0;
   end else begin
       if ((dat_rsp_exec_pvld_d5) == 1'b1) begin
           dat_rsp_exec_dummy_d6 <= dat_rsp_exec_dummy_d5;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d5) == 1'b0) begin
       end else begin
           dat_rsp_exec_dummy_d6 <= 'bx;
       // VCS coverage on
       end
   end
end
reg [1:0] dat_rsp_exec_sub_h_d6;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_exec_sub_h_d6 <= {2{1'b0}};
   end else begin
       if ((dat_rsp_exec_pvld_d5) == 1'b1) begin
           dat_rsp_exec_sub_h_d6 <= dat_rsp_exec_sub_h_d5;
       // VCS coverage off
       end else if ((dat_rsp_exec_pvld_d5) == 1'b0) begin
       end else begin
           dat_rsp_exec_sub_h_d6 <= 'bx;
       // VCS coverage on
       end
   end
end
assign dat_rsp_pipe_pvld = dat_rsp_pipe_pvld_d6;
assign dat_rsp_pipe_pd = dat_rsp_pipe_pd_d6;
assign dat_rsp_exec_pvld = dat_rsp_exec_pvld_d6;
assign dat_rsp_exec_dummy = dat_rsp_exec_dummy_d6;
assign dat_rsp_exec_sub_h = dat_rsp_exec_sub_h_d6;


//| eperl: generated_end (DO NOT EDIT ABOVE)
// PKT_UNPACK_WIRE( csc_dat_req_pkg , dat_rsp_pipe_ , dat_rsp_pipe_pd )
assign dat_rsp_pipe_sub_w[1:0] = dat_rsp_pipe_pd[1:0];
assign dat_rsp_pipe_sub_h[1:0] = dat_rsp_pipe_pd[3:2];
assign dat_rsp_pipe_sub_c = dat_rsp_pipe_pd[4];
assign dat_rsp_pipe_ch_end = dat_rsp_pipe_pd[5];
assign dat_rsp_pipe_bytes[7:0] = dat_rsp_pipe_pd[14:7];
assign dat_rsp_pipe_cur_sub_h[1:0] = dat_rsp_pipe_pd[16:15];
assign dat_rsp_pipe_dummy = dat_rsp_pipe_pd[17];
assign dat_rsp_pipe_sub_w_st = dat_rsp_pipe_pd[18];
assign dat_rsp_pipe_rls = dat_rsp_pipe_pd[19];
assign dat_rsp_pipe_flag[8:0] = dat_rsp_pipe_pd[28:20];
//////////////////////////////////////////////////////////////
///// dl data cache                                      /////
//////////////////////////////////////////////////////////////
assign dat_l0c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h0));
assign dat_l1c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h1));
assign dat_l2c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h2));
assign dat_l3c0_en = (sc2buf_dat_rd_valid & (dat_rsp_exec_sub_h == 2'h3));
//only winograd/image
assign dat_l0c1_en = (dat_wg_adv & ~dat_rsp_exec_sub_h[0]) | (is_img_d1[12] & dat_l0c0_en & ~dat_l0c0_dummy);
assign dat_l1c1_en = (dat_wg_adv & dat_rsp_exec_sub_h[0]) | (is_img_d1[13] & dat_l1c0_en & ~dat_l1c0_dummy);
assign dat_l2c1_en = (is_img_d1[15] & dat_l2c0_en & ~dat_l2c0_dummy);
assign dat_l3c1_en = (is_img_d1[16] & dat_l3c0_en & ~dat_l3c0_dummy);
assign dat_dummy_l0_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h0);
assign dat_dummy_l1_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h1);
assign dat_dummy_l2_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h2);
assign dat_dummy_l3_en = dat_rsp_exec_pvld & dat_rsp_exec_dummy & (dat_rsp_exec_sub_h == 2'h3);
assign dat_wg_adv = sc2buf_dat_rd_valid & is_winograd_d1[11] & ~dat_rsp_pipe_sub_w_st;
assign dat_l0c0_dummy_w = dat_l0c0_en ? 1'b0 : dat_dummy_l0_en ? 1'b1 : dat_l0c0_dummy;
assign dat_l1c0_dummy_w = dat_l1c0_en ? 1'b0 : dat_dummy_l1_en ? 1'b1 : dat_l1c0_dummy;
assign dat_l2c0_dummy_w = dat_l2c0_en ? 1'b0 : dat_dummy_l2_en ? 1'b1 : dat_l2c0_dummy;
assign dat_l3c0_dummy_w = dat_l3c0_en ? 1'b0 : dat_dummy_l3_en ? 1'b1 : dat_l3c0_dummy;
assign dat_l0c1_dummy_w = dat_l0c1_en ? 1'b0 : (dat_l0_set) ? dat_l0c0_dummy : dat_l0c1_dummy;
assign dat_l1c1_dummy_w = dat_l1c1_en ? 1'b0 : (dat_l1_set & (|sub_h_total_g2)) ? dat_l1c0_dummy : dat_l1c1_dummy;
assign dat_l2c1_dummy_w = dat_l2c1_en ? 1'b0 : (dat_l2_set & sub_h_total_g2[1]) ? dat_l2c0_dummy : dat_l2c1_dummy;
assign dat_l3c1_dummy_w = dat_l3c1_en ? 1'b0 : (dat_l3_set & sub_h_total_g2[1]) ? dat_l3c0_dummy : dat_l3c1_dummy;
assign dat_l0_set = dat_l0c0_en | dat_dummy_l0_en;
assign dat_l1_set = dat_l1c0_en | dat_dummy_l1_en;
assign dat_l2_set = dat_l2c0_en | dat_dummy_l2_en;
assign dat_l3_set = dat_l3c0_en | dat_dummy_l3_en;
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l0c0_dummy_w\" -q dat_l0c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l1c0_dummy_w\" -q dat_l1c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l2c0_dummy_w\" -q dat_l2c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l3c0_dummy_w\" -q dat_l3c0_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l0c1_dummy_w\" -q dat_l0c1_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l1c1_dummy_w\" -q dat_l1c1_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l2c1_dummy_w\" -q dat_l2c1_dummy");
//: &eperl::flop("-nodeclare   -rval \"1'b1\"   -d \"dat_l3c1_dummy_w\" -q dat_l3c1_dummy");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l0c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l0c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l1c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l1c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l2c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l2c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l3c0_en\" -d \"sc2buf_dat_rd_data\" -q dat_l3c0 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l0c1_en\" -d dat_l0c0 -q dat_l0c1 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l1c1_en\" -d dat_l1c0 -q dat_l1c1 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l2c1_en\" -d dat_l2c0 -q dat_l2c1 ");
//: &eperl::flop("-nodeclare  -norst -en \"dat_l3c1_en\" -d dat_l3c0 -q dat_l3c1 ");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l0c0_dummy <= 1'b1;
   end else begin
       dat_l0c0_dummy <= dat_l0c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l1c0_dummy <= 1'b1;
   end else begin
       dat_l1c0_dummy <= dat_l1c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l2c0_dummy <= 1'b1;
   end else begin
       dat_l2c0_dummy <= dat_l2c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l3c0_dummy <= 1'b1;
   end else begin
       dat_l3c0_dummy <= dat_l3c0_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l0c1_dummy <= 1'b1;
   end else begin
       dat_l0c1_dummy <= dat_l0c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l1c1_dummy <= 1'b1;
   end else begin
       dat_l1c1_dummy <= dat_l1c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l2c1_dummy <= 1'b1;
   end else begin
       dat_l2c1_dummy <= dat_l2c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_l3c1_dummy <= 1'b1;
   end else begin
       dat_l3c1_dummy <= dat_l3c1_dummy_w;
   end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l0c0_en) == 1'b1) begin
           dat_l0c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l0c0_en) == 1'b0) begin
       end else begin
           dat_l0c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l1c0_en) == 1'b1) begin
           dat_l1c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l1c0_en) == 1'b0) begin
       end else begin
           dat_l1c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l2c0_en) == 1'b1) begin
           dat_l2c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l2c0_en) == 1'b0) begin
       end else begin
           dat_l2c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l3c0_en) == 1'b1) begin
           dat_l3c0 <= sc2buf_dat_rd_data;
       // VCS coverage off
       end else if ((dat_l3c0_en) == 1'b0) begin
       end else begin
           dat_l3c0 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l0c1_en) == 1'b1) begin
           dat_l0c1 <= dat_l0c0;
       // VCS coverage off
       end else if ((dat_l0c1_en) == 1'b0) begin
       end else begin
           dat_l0c1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l1c1_en) == 1'b1) begin
           dat_l1c1 <= dat_l1c0;
       // VCS coverage off
       end else if ((dat_l1c1_en) == 1'b0) begin
       end else begin
           dat_l1c1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l2c1_en) == 1'b1) begin
           dat_l2c1 <= dat_l2c0;
       // VCS coverage off
       end else if ((dat_l2c1_en) == 1'b0) begin
       end else begin
           dat_l2c1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_l3c1_en) == 1'b1) begin
           dat_l3c1 <= dat_l3c0;
       // VCS coverage off
       end else if ((dat_l3c1_en) == 1'b0) begin
       end else begin
           dat_l3c1 <= 'bx;
       // VCS coverage on
       end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// response contorl                                   /////
//////////////////////////////////////////////////////////////
// PKT_PACK_WIRE( csc_dat_rsp_pkg , dat_rsp_pipe_ , dat_rsp_pd_d0 )
assign dat_rsp_pd_d0[1:0] = dat_rsp_pipe_sub_w[1:0];
assign dat_rsp_pd_d0[3:2] = dat_rsp_pipe_sub_h[1:0];
assign dat_rsp_pd_d0[4] = dat_rsp_pipe_sub_c ;
assign dat_rsp_pd_d0[5] = dat_rsp_pipe_ch_end ;
assign dat_rsp_pd_d0[6] = 1'b0 ;
assign dat_rsp_pd_d0[14:7] = dat_rsp_pipe_bytes[7:0];
assign dat_rsp_pd_d0[16:15] = dat_rsp_pipe_cur_sub_h[1:0];
assign dat_rsp_pd_d0[17] = dat_rsp_pipe_rls ;
assign dat_rsp_pd_d0[26:18] = dat_rsp_pipe_flag[8:0];
//add latency
//: my $delay_depth = 4;
//: my $i;
//: my $j;
//:
//: print "assign dat_rsp_pvld_d0 = dat_rsp_pipe_pvld;\n";
//: for($i = 0; $i < $delay_depth; $i ++) {
//: $j = $i + 1;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"           -d \"dat_rsp_pvld_d${i}\"   -q dat_rsp_pvld_d${j}");
//: &eperl::flop("-nodeclare   -rval \"{27{1'b0}}\"     -en \"dat_rsp_pvld_d${i}\"  -d \"dat_rsp_pd_d${i}\" -q dat_rsp_pd_d${j}");
//: }
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_rsp_pvld_d0 = dat_rsp_pipe_pvld;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d1 <= 1'b0;
   end else begin
       dat_rsp_pvld_d1 <= dat_rsp_pvld_d0;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d1 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d0) == 1'b1) begin
           dat_rsp_pd_d1 <= dat_rsp_pd_d0;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d0) == 1'b0) begin
       end else begin
           dat_rsp_pd_d1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d2 <= 1'b0;
   end else begin
       dat_rsp_pvld_d2 <= dat_rsp_pvld_d1;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d2 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d1) == 1'b1) begin
           dat_rsp_pd_d2 <= dat_rsp_pd_d1;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d1) == 1'b0) begin
       end else begin
           dat_rsp_pd_d2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d3 <= 1'b0;
   end else begin
       dat_rsp_pvld_d3 <= dat_rsp_pvld_d2;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d3 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d2) == 1'b1) begin
           dat_rsp_pd_d3 <= dat_rsp_pd_d2;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d2) == 1'b0) begin
       end else begin
           dat_rsp_pd_d3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pvld_d4 <= 1'b0;
   end else begin
       dat_rsp_pvld_d4 <= dat_rsp_pvld_d3;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_rsp_pd_d4 <= {27{1'b0}};
   end else begin
       if ((dat_rsp_pvld_d3) == 1'b1) begin
           dat_rsp_pd_d4 <= dat_rsp_pd_d3;
       // VCS coverage off
       end else if ((dat_rsp_pvld_d3) == 1'b0) begin
       end else begin
           dat_rsp_pd_d4 <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dat_rsp_pvld = (sub_h_total_g3[2] & dat_rsp_pvld_d4) |
                      (sub_h_total_g3[1] & dat_rsp_pvld_d2) |
                      (sub_h_total_g3[0] & dat_rsp_pvld_d1);
assign dat_rsp_l0_pvld = dat_rsp_pvld_d1;
assign dat_rsp_l1_pvld = dat_rsp_pvld_d2;
assign dat_rsp_l2_pvld = dat_rsp_pvld_d3;
assign dat_rsp_l3_pvld = dat_rsp_pvld_d4;
assign dat_rsp_pd = ({27 {sub_h_total_g4[2]}} & dat_rsp_pd_d4) |
                    ({27 {sub_h_total_g4[1]}} & dat_rsp_pd_d2) |
                    ({27 {sub_h_total_g4[0]}} & dat_rsp_pd_d1);
assign dat_rsp_l0_sub_c = dat_rsp_pd_d1[4:4];
assign dat_rsp_l1_sub_c = dat_rsp_pd_d2[4:4];
assign dat_rsp_l2_sub_c = dat_rsp_pd_d3[4:4];
assign dat_rsp_l3_sub_c = dat_rsp_pd_d4[4:4];
assign dat_rsp_l0_flag = dat_rsp_pd_d1[26:18];
assign dat_rsp_l1_flag = dat_rsp_pd_d2[26:18];
assign dat_rsp_l2_flag = dat_rsp_pd_d3[26:18];
assign dat_rsp_l3_flag = dat_rsp_pd_d4[26:18];
assign dat_rsp_l0_stripe_end = dat_rsp_l0_flag[6:6];
assign dat_rsp_l1_stripe_end = dat_rsp_l1_flag[6:6];
assign dat_rsp_l2_stripe_end = dat_rsp_l2_flag[6:6];
assign dat_rsp_l3_stripe_end = dat_rsp_l3_flag[6:6];
// PKT_UNPACK_WIRE( csc_dat_rsp_pkg , dat_rsp_ , dat_rsp_pd )
assign dat_rsp_sub_w[1:0] = dat_rsp_pd[1:0];
assign dat_rsp_sub_h[1:0] = dat_rsp_pd[3:2];
assign dat_rsp_sub_c = dat_rsp_pd[4];
assign dat_rsp_ch_end = dat_rsp_pd[5];
assign dat_rsp_bytes[7:0] = dat_rsp_pd[14:7];
assign dat_rsp_cur_sub_h[1:0] = dat_rsp_pd[16:15];
assign dat_rsp_rls = dat_rsp_pd[17];
assign dat_rsp_flag[8:0] = dat_rsp_pd[26:18];
// PKT_UNPACK_WIRE( nvdla_stripe_info , dat_rsp_ , dat_rsp_flag )
assign dat_rsp_batch_index[4:0] = dat_rsp_flag[4:0];
assign dat_rsp_stripe_st = dat_rsp_flag[5];
assign dat_rsp_stripe_end = dat_rsp_flag[6];
assign dat_rsp_channel_end = dat_rsp_flag[7];
assign dat_rsp_layer_end = dat_rsp_flag[8];
assign rsp_sft_cnt_l0_sub = dat_l0c0_en ? 8'h40   : 8'h0;
assign rsp_sft_cnt_l1_sub = dat_l1c0_en ? 8'h40   : 8'h0;
assign rsp_sft_cnt_l2_sub = dat_l2c0_en ? 8'h40   : 8'h0;
assign rsp_sft_cnt_l3_sub = dat_l3c0_en ? 8'h40   : 8'h0;
////: &eperl::retime("-O stripe_begin_disable_jump_7T -i stripe_begin_disable_jump -stage 8 -clk nvdla_core_clk");
////: &eperl::flop("-q stripe_begin_disable_jump_8T -d stripe_begin_disable_jump_7T -clk nvdla_core_clk");
assign {mon_rsp_sft_cnt_l0_w,rsp_sft_cnt_l0_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l0 + pixel_x_byte_stride - rsp_sft_cnt_l0_sub);
assign {mon_rsp_sft_cnt_l1_w,rsp_sft_cnt_l1_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l1 + pixel_x_byte_stride - rsp_sft_cnt_l1_sub);
assign {mon_rsp_sft_cnt_l2_w,rsp_sft_cnt_l2_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l2 + pixel_x_byte_stride - rsp_sft_cnt_l2_sub);
assign {mon_rsp_sft_cnt_l3_w,rsp_sft_cnt_l3_inc} = (pixel_x_byte_stride > 8'h40  ) ? 8'h40   :
                                                    (rsp_sft_cnt_l3 + pixel_x_byte_stride - rsp_sft_cnt_l3_sub);
//the data frm cbuf's low Bytes is always needed. High Bytes maybe unneeded.
assign dat_rsp_l0_block_end = dat_rsp_l0_sub_c;
assign dat_rsp_l1_block_end = dat_rsp_l1_sub_c;
assign dat_rsp_l2_block_end = dat_rsp_l2_sub_c;
assign dat_rsp_l3_block_end = dat_rsp_l3_sub_c;
assign rsp_sft_cnt_l0_w = (layer_st) ? 8'h40   : //begin from C0
                          (dat_rsp_l0_stripe_end & ~dat_rsp_l0_block_end) ? rsp_sft_cnt_l0_ori :
                          (dat_rsp_l0_stripe_end & dat_rsp_l0_block_end) ? 8'h40   :
                          (dat_dummy_l0_en) ? (rsp_sft_cnt_l0_inc & 8'h3f) :
                          rsp_sft_cnt_l0_inc;
assign rsp_sft_cnt_l1_w = (layer_st) ? 8'h40   :
                          (dat_rsp_l1_stripe_end & ~dat_rsp_l1_block_end) ? rsp_sft_cnt_l1_ori :
                          (dat_rsp_l1_stripe_end & dat_rsp_l1_block_end) ? 8'h40   :
                          (dat_dummy_l1_en) ? (rsp_sft_cnt_l1_inc & 8'h3f) :
                          rsp_sft_cnt_l1_inc;
assign rsp_sft_cnt_l2_w = (layer_st) ? 8'h40   :
                          (dat_rsp_l2_stripe_end & ~dat_rsp_l2_block_end) ? rsp_sft_cnt_l2_ori :
                          (dat_rsp_l2_stripe_end & dat_rsp_l2_block_end) ? 8'h40   :
                          (dat_dummy_l2_en) ? (rsp_sft_cnt_l2_inc & 8'h3f) :
                          rsp_sft_cnt_l2_inc;
assign rsp_sft_cnt_l3_w = (layer_st) ? 8'h40   :
                          (dat_rsp_l3_stripe_end & ~dat_rsp_l3_block_end) ? rsp_sft_cnt_l3_ori :
                          (dat_rsp_l3_stripe_end & dat_rsp_l3_block_end) ? 8'h40   :
                          (dat_dummy_l3_en) ? (rsp_sft_cnt_l3_inc & 8'h3f) :
                          rsp_sft_cnt_l3_inc;
assign rsp_sft_cnt_l0_en = layer_st | (is_img_d1[17] & dat_rsp_l0_pvld);
assign rsp_sft_cnt_l1_en = layer_st | (is_img_d1[18] & dat_rsp_l1_pvld & (sub_h_total_g5 != 3'h1));
assign rsp_sft_cnt_l2_en = layer_st | (is_img_d1[19] & dat_rsp_l2_pvld & (sub_h_total_g5 == 3'h4));
assign rsp_sft_cnt_l3_en = layer_st | (is_img_d1[20] & dat_rsp_l3_pvld & (sub_h_total_g5 == 3'h4));
assign rsp_sft_cnt_l0_ori_en = layer_st | (is_img_d1[21] & dat_rsp_l0_pvld & dat_rsp_l0_stripe_end & dat_rsp_l0_block_end);
assign rsp_sft_cnt_l1_ori_en = layer_st | (is_img_d1[22] & dat_rsp_l1_pvld & dat_rsp_l1_stripe_end & dat_rsp_l1_block_end & (sub_h_total_g6 != 3'h1));
assign rsp_sft_cnt_l2_ori_en = layer_st | (is_img_d1[23] & dat_rsp_l2_pvld & dat_rsp_l2_stripe_end & dat_rsp_l2_block_end & (sub_h_total_g6 == 3'h4));
assign rsp_sft_cnt_l3_ori_en = layer_st | (is_img_d1[24] & dat_rsp_l3_pvld & dat_rsp_l3_stripe_end & dat_rsp_l3_block_end & (sub_h_total_g6 == 3'h4));
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l0_en\" -d \"rsp_sft_cnt_l0_w\" -q rsp_sft_cnt_l0");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l1_en\" -d \"rsp_sft_cnt_l1_w\" -q rsp_sft_cnt_l1");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l2_en\" -d \"rsp_sft_cnt_l2_w\" -q rsp_sft_cnt_l2");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l3_en\" -d \"rsp_sft_cnt_l3_w\" -q rsp_sft_cnt_l3");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l0_ori_en\" -d \"rsp_sft_cnt_l0_w\" -q rsp_sft_cnt_l0_ori");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l1_ori_en\" -d \"rsp_sft_cnt_l1_w\" -q rsp_sft_cnt_l1_ori");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l2_ori_en\" -d \"rsp_sft_cnt_l2_w\" -q rsp_sft_cnt_l2_ori");
//: &eperl::flop("-nodeclare   -rval \"{8{1'b0}}\"  -en \"rsp_sft_cnt_l3_ori_en\" -d \"rsp_sft_cnt_l3_w\" -q rsp_sft_cnt_l3_ori");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l0 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l0_en) == 1'b1) begin
           rsp_sft_cnt_l0 <= rsp_sft_cnt_l0_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l0_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l0 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l1 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l1_en) == 1'b1) begin
           rsp_sft_cnt_l1 <= rsp_sft_cnt_l1_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l1_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l1 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l2 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l2_en) == 1'b1) begin
           rsp_sft_cnt_l2 <= rsp_sft_cnt_l2_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l2_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l2 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l3 <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l3_en) == 1'b1) begin
           rsp_sft_cnt_l3 <= rsp_sft_cnt_l3_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l3_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l3 <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l0_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l0_ori_en) == 1'b1) begin
           rsp_sft_cnt_l0_ori <= rsp_sft_cnt_l0_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l0_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l0_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l1_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l1_ori_en) == 1'b1) begin
           rsp_sft_cnt_l1_ori <= rsp_sft_cnt_l1_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l1_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l1_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l2_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l2_ori_en) == 1'b1) begin
           rsp_sft_cnt_l2_ori <= rsp_sft_cnt_l2_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l2_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l2_ori <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       rsp_sft_cnt_l3_ori <= {8{1'b0}};
   end else begin
       if ((rsp_sft_cnt_l3_ori_en) == 1'b1) begin
           rsp_sft_cnt_l3_ori <= rsp_sft_cnt_l3_w;
       // VCS coverage off
       end else if ((rsp_sft_cnt_l3_ori_en) == 1'b0) begin
       end else begin
           rsp_sft_cnt_l3_ori <= 'bx;
       // VCS coverage on
       end
   end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// response data                                      /////
//////////////////////////////////////////////////////////////
//////////////// data for winograd ////////////////
//winograd need future update

//////////////// data for convlution ////////////////
assign dat_rsp_pad_value = {64{pad_value[7:0]}};
assign dat_rsp_l0c0 = dat_l0c0_dummy ? dat_rsp_pad_value : dat_l0c0;
assign dat_rsp_l1c0 = dat_l1c0_dummy ? dat_rsp_pad_value : dat_l1c0;
assign dat_rsp_l2c0 = dat_l2c0_dummy ? dat_rsp_pad_value : dat_l2c0;
assign dat_rsp_l3c0 = dat_l3c0_dummy ? dat_rsp_pad_value : dat_l3c0;
assign dat_rsp_l0c1 = dat_l0c1_dummy ? dat_rsp_pad_value : dat_l0c1;
assign dat_rsp_l1c1 = dat_l1c1_dummy ? dat_rsp_pad_value : dat_l1c1;
assign dat_rsp_l2c1 = dat_l2c1_dummy ? dat_rsp_pad_value : dat_l2c1;
assign dat_rsp_l3c1 = dat_l3c1_dummy ? dat_rsp_pad_value : dat_l3c1;
//several atomM may combine together as an entry

assign dat_rsp_conv_8b = (is_winograd_d1[14] | is_img_d1[26]) ? {512{1'b0}} :
((dat_rsp_bytes <= 8'h20)&((dat_rsp_sub_w[0] == 1'h0))) ? {{512/2{1'b0}}, dat_rsp_l0c0[512/2 -1:0]} :
((dat_rsp_bytes <= 8'h20)&((dat_rsp_sub_w[0] == 1'h1))) ? {{512/2{1'b0}}, dat_rsp_l0c0[512 -1:512/2]} :
                dat_rsp_l0c0;
assign dat_rsp_conv = dat_rsp_conv_8b;
//////////////// data for image ////////////////
assign dat_rsp_l0_sft_in = ~is_img_d1[27] ? 'b0 : {dat_rsp_l0c0, dat_rsp_l0c1};
assign dat_rsp_l1_sft_in = ~is_img_d1[28] ? 'b0 : {dat_rsp_l1c0, dat_rsp_l1c1};
assign dat_rsp_l2_sft_in = ~is_img_d1[29] ? 'b0 : {dat_rsp_l2c0, dat_rsp_l2c1};
assign dat_rsp_l3_sft_in = ~is_img_d1[30] ? 'b0 : {dat_rsp_l3c0, dat_rsp_l3c1};
assign {mon_dat_rsp_l0_sft, dat_rsp_l0_sft} = dat_rsp_l0_sft_in >> {rsp_sft_cnt_l0, 3'b0};
assign {mon_dat_rsp_l1_sft, dat_rsp_l1_sft} = dat_rsp_l1_sft_in >> {rsp_sft_cnt_l1, 3'b0};
assign {mon_dat_rsp_l2_sft, dat_rsp_l2_sft} = dat_rsp_l2_sft_in >> {rsp_sft_cnt_l2, 3'b0};
assign {mon_dat_rsp_l3_sft, dat_rsp_l3_sft} = dat_rsp_l3_sft_in >> {rsp_sft_cnt_l3, 3'b0};
assign dat_rsp_img_8b = (~is_img_d1[32])? 'b0 :
                        (sub_h_total_g8 == 3'h4) ? {dat_rsp_l3_sft[512/4 -1:0], dat_rsp_l2_sft_d3[512/4 -1:0], dat_rsp_l1_sft_d3[512/4 -1:0], dat_rsp_l0_sft_d3[512/4 -1:0]} :
                        (sub_h_total_g8 == 3'h2) ? {dat_rsp_l1_sft[512/2 -1:0], dat_rsp_l0_sft_d1[512/2 -1:0]} :
                        dat_rsp_l0_sft[512 -1:0];
assign dat_rsp_img = dat_rsp_img_8b;
wire dat_rsp_sft_d1_en = dat_rsp_l0_pvld & (sub_h_total_g9 != 3'h1);
wire dat_rsp_sft_d2_en = dat_rsp_l1_pvld & (sub_h_total_g9 == 3'h4);
wire dat_rsp_sft_d3_en = dat_rsp_l2_pvld & (sub_h_total_g9 == 3'h4);
//: my $half=512/2;
//: my $quat=512/4;
//: &eperl::flop("-nodeclare -wid ${half} -norst -en \"dat_rsp_sft_d1_en\" -d \"dat_rsp_l0_sft\" -q dat_rsp_l0_sft_d1");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d2_en\" -d \"dat_rsp_l0_sft_d1\" -q dat_rsp_l0_sft_d2");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d3_en\" -d \"dat_rsp_l0_sft_d2\" -q dat_rsp_l0_sft_d3");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d2_en\" -d \"dat_rsp_l1_sft\" -q dat_rsp_l1_sft_d2");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d3_en\" -d \"dat_rsp_l1_sft_d2\" -q dat_rsp_l1_sft_d3");
//: &eperl::flop("-nodeclare -wid ${quat} -norst -en \"dat_rsp_sft_d3_en\" -d \"dat_rsp_l2_sft\" -q dat_rsp_l2_sft_d3");
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d1_en) == 1'b1) begin
           dat_rsp_l0_sft_d1 <= dat_rsp_l0_sft;
       // VCS coverage off
       end else if ((dat_rsp_sft_d1_en) == 1'b0) begin
       end else begin
           dat_rsp_l0_sft_d1 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d2_en) == 1'b1) begin
           dat_rsp_l0_sft_d2 <= dat_rsp_l0_sft_d1;
       // VCS coverage off
       end else if ((dat_rsp_sft_d2_en) == 1'b0) begin
       end else begin
           dat_rsp_l0_sft_d2 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d3_en) == 1'b1) begin
           dat_rsp_l0_sft_d3 <= dat_rsp_l0_sft_d2;
       // VCS coverage off
       end else if ((dat_rsp_sft_d3_en) == 1'b0) begin
       end else begin
           dat_rsp_l0_sft_d3 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d2_en) == 1'b1) begin
           dat_rsp_l1_sft_d2 <= dat_rsp_l1_sft;
       // VCS coverage off
       end else if ((dat_rsp_sft_d2_en) == 1'b0) begin
       end else begin
           dat_rsp_l1_sft_d2 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d3_en) == 1'b1) begin
           dat_rsp_l1_sft_d3 <= dat_rsp_l1_sft_d2;
       // VCS coverage off
       end else if ((dat_rsp_sft_d3_en) == 1'b0) begin
       end else begin
           dat_rsp_l1_sft_d3 <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_rsp_sft_d3_en) == 1'b1) begin
           dat_rsp_l2_sft_d3 <= dat_rsp_l2_sft;
       // VCS coverage off
       end else if ((dat_rsp_sft_d3_en) == 1'b0) begin
       end else begin
           dat_rsp_l2_sft_d3 <= 'bx;
       // VCS coverage on
       end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////// byte mask ////////////////
//sub_h_total=2, each sub_h align to 1/2 entry;
//sub_h_total=4, each sub_h align to 1/4 entry;
assign dat_rsp_ori_mask = ~({64{1'b1}} << dat_rsp_bytes);
assign dat_rsp_cur_h_mask_p1 = (dat_rsp_cur_sub_h >= 2'h1) ? {64{1'b1}} : 'b0;
assign dat_rsp_cur_h_mask_p2 = (dat_rsp_cur_sub_h >= 2'h2) ? {64/2{1'b1}} : 'b0;
assign dat_rsp_cur_h_mask_p3 = (dat_rsp_cur_sub_h == 2'h3) ? {64/2{1'b1}} : 'b0;
assign dat_rsp_cur_h_e2_mask_8b = {dat_rsp_cur_h_mask_p1[64/2 -1:0], {64/2{1'b1}}};
assign dat_rsp_cur_h_e4_mask_8b = {dat_rsp_cur_h_mask_p3[64/4 -1:0], dat_rsp_cur_h_mask_p2[64/4 -1:0], dat_rsp_cur_h_mask_p1[64/4 -1:0], {64/4{1'b1}}};
assign dat_rsp_mask_8b = (sub_h_total_g11 == 3'h4) ? ({4{dat_rsp_ori_mask[64/4 -1:0]}} & dat_rsp_cur_h_e4_mask_8b) :
                         (sub_h_total_g11 == 3'h2) ? ({2{dat_rsp_ori_mask[64/2 -1:0]}} & dat_rsp_cur_h_e2_mask_8b) :
                         dat_rsp_ori_mask[64 -1:0];
assign dat_rsp_data_w = is_img_d1[33] ? dat_rsp_img :
                        dat_rsp_conv;
//: my $i;
//: my $b1;
//: my $b0;
//: my $kk=64 -1;
//: print "assign dat_rsp_mask_val_int8 = {";
//: for($i = ${kk}; $i >= 0; $i --) {
//: $b0 = sprintf("%3d", $i * 8);
//: $b1 = sprintf("%3d", $i * 8 + 7);
//: print "(|dat_rsp_data_w[${b1}:${b0}])";
//: if($i == 0) {
//: print "};\n";
//: } elsif ($i % 8 == 0) {
//: print ",\n                               ";
//: } else {
//: print ", ";
//: }
//: }
//: print "\n\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_rsp_mask_val_int8 = {(|dat_rsp_data_w[511:504]), (|dat_rsp_data_w[503:496]), (|dat_rsp_data_w[495:488]), (|dat_rsp_data_w[487:480]), (|dat_rsp_data_w[479:472]), (|dat_rsp_data_w[471:464]), (|dat_rsp_data_w[463:456]), (|dat_rsp_data_w[455:448]),
                               (|dat_rsp_data_w[447:440]), (|dat_rsp_data_w[439:432]), (|dat_rsp_data_w[431:424]), (|dat_rsp_data_w[423:416]), (|dat_rsp_data_w[415:408]), (|dat_rsp_data_w[407:400]), (|dat_rsp_data_w[399:392]), (|dat_rsp_data_w[391:384]),
                               (|dat_rsp_data_w[383:376]), (|dat_rsp_data_w[375:368]), (|dat_rsp_data_w[367:360]), (|dat_rsp_data_w[359:352]), (|dat_rsp_data_w[351:344]), (|dat_rsp_data_w[343:336]), (|dat_rsp_data_w[335:328]), (|dat_rsp_data_w[327:320]),
                               (|dat_rsp_data_w[319:312]), (|dat_rsp_data_w[311:304]), (|dat_rsp_data_w[303:296]), (|dat_rsp_data_w[295:288]), (|dat_rsp_data_w[287:280]), (|dat_rsp_data_w[279:272]), (|dat_rsp_data_w[271:264]), (|dat_rsp_data_w[263:256]),
                               (|dat_rsp_data_w[255:248]), (|dat_rsp_data_w[247:240]), (|dat_rsp_data_w[239:232]), (|dat_rsp_data_w[231:224]), (|dat_rsp_data_w[223:216]), (|dat_rsp_data_w[215:208]), (|dat_rsp_data_w[207:200]), (|dat_rsp_data_w[199:192]),
                               (|dat_rsp_data_w[191:184]), (|dat_rsp_data_w[183:176]), (|dat_rsp_data_w[175:168]), (|dat_rsp_data_w[167:160]), (|dat_rsp_data_w[159:152]), (|dat_rsp_data_w[151:144]), (|dat_rsp_data_w[143:136]), (|dat_rsp_data_w[135:128]),
                               (|dat_rsp_data_w[127:120]), (|dat_rsp_data_w[119:112]), (|dat_rsp_data_w[111:104]), (|dat_rsp_data_w[103: 96]), (|dat_rsp_data_w[ 95: 88]), (|dat_rsp_data_w[ 87: 80]), (|dat_rsp_data_w[ 79: 72]), (|dat_rsp_data_w[ 71: 64]),
                               (|dat_rsp_data_w[ 63: 56]), (|dat_rsp_data_w[ 55: 48]), (|dat_rsp_data_w[ 47: 40]), (|dat_rsp_data_w[ 39: 32]), (|dat_rsp_data_w[ 31: 24]), (|dat_rsp_data_w[ 23: 16]), (|dat_rsp_data_w[ 15:  8]), (|dat_rsp_data_w[  7:  0])};



//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dat_rsp_mask_w = (dat_rsp_mask_8b & dat_rsp_mask_val_int8) ;
assign dat_rsp_p1_vld_w = 1'b0;
assign dat_rsp_p0_vld_w = dat_rsp_pvld & ~is_winograd_d1[16];
//////////////////////////////////////////////////////////////
///// latency register to balance with PRA cell          /////
//////////////////////////////////////////////////////////////
//: my $total_latency = 5;
//:
//: print "assign dat_out_pvld_l0 = dat_rsp_pvld;\n";
//: print "assign dat_out_flag_l0 = dat_rsp_flag;\n";
//: for(my $i = 0; $i < $total_latency; $i ++) {
//: my $j = $i + 1;
//: &eperl::flop("-wid 1   -rval \"1'b0\"       -d \"dat_out_pvld_l${i}\"   -q dat_out_pvld_l${j}");
//: &eperl::flop("-wid 9   -rval \"{9{1'b0}}\"  -en \"dat_out_pvld_l${i}\"  -d \"dat_out_flag_l${i}\" -q dat_out_flag_l${j}");
//: }
//:
//: my $k = $total_latency;
//: print "assign dat_out_pvld_w = is_winograd_d1[17] ? dat_out_pvld_l${k} : dat_rsp_pvld;\n";
//: print "assign dat_out_flag_w = is_winograd_d1[18] ? dat_out_flag_l${k} : dat_rsp_flag;\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
assign dat_out_pvld_l0 = dat_rsp_pvld;
assign dat_out_flag_l0 = dat_rsp_flag;
reg  dat_out_pvld_l1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l1 <= 1'b0;
   end else begin
       dat_out_pvld_l1 <= dat_out_pvld_l0;
   end
end
reg [8:0] dat_out_flag_l1;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l1 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l0) == 1'b1) begin
           dat_out_flag_l1 <= dat_out_flag_l0;
       // VCS coverage off
       end else if ((dat_out_pvld_l0) == 1'b0) begin
       end else begin
           dat_out_flag_l1 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l2 <= 1'b0;
   end else begin
       dat_out_pvld_l2 <= dat_out_pvld_l1;
   end
end
reg [8:0] dat_out_flag_l2;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l2 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l1) == 1'b1) begin
           dat_out_flag_l2 <= dat_out_flag_l1;
       // VCS coverage off
       end else if ((dat_out_pvld_l1) == 1'b0) begin
       end else begin
           dat_out_flag_l2 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l3 <= 1'b0;
   end else begin
       dat_out_pvld_l3 <= dat_out_pvld_l2;
   end
end
reg [8:0] dat_out_flag_l3;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l3 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l2) == 1'b1) begin
           dat_out_flag_l3 <= dat_out_flag_l2;
       // VCS coverage off
       end else if ((dat_out_pvld_l2) == 1'b0) begin
       end else begin
           dat_out_flag_l3 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l4 <= 1'b0;
   end else begin
       dat_out_pvld_l4 <= dat_out_pvld_l3;
   end
end
reg [8:0] dat_out_flag_l4;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l4 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l3) == 1'b1) begin
           dat_out_flag_l4 <= dat_out_flag_l3;
       // VCS coverage off
       end else if ((dat_out_pvld_l3) == 1'b0) begin
       end else begin
           dat_out_flag_l4 <= 'bx;
       // VCS coverage on
       end
   end
end
reg  dat_out_pvld_l5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld_l5 <= 1'b0;
   end else begin
       dat_out_pvld_l5 <= dat_out_pvld_l4;
   end
end
reg [8:0] dat_out_flag_l5;
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag_l5 <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_l4) == 1'b1) begin
           dat_out_flag_l5 <= dat_out_flag_l4;
       // VCS coverage off
       end else if ((dat_out_pvld_l4) == 1'b0) begin
       end else begin
           dat_out_flag_l5 <= 'bx;
       // VCS coverage on
       end
   end
end
assign dat_out_pvld_w = is_winograd_d1[17] ? dat_out_pvld_l5 : dat_rsp_pvld;
assign dat_out_flag_w = is_winograd_d1[18] ? dat_out_flag_l5 : dat_rsp_flag;

//| eperl: generated_end (DO NOT EDIT ABOVE)
assign dat_out_bypass_p0_vld_w = dat_rsp_p0_vld_w;
assign dat_out_bypass_mask_w = dat_rsp_mask_w;
assign dat_out_bypass_data_w = dat_rsp_data_w;
//: my $kk=64;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_out_pvld_w\" -q dat_out_pvld");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_out_pvld_w\" -d \"dat_out_flag_w\" -q dat_out_flag");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dat_out_bypass_p0_vld_w\" -d \"dat_out_bypass_mask_w\" -q dat_out_bypass_mask");
//: for(my $i = 0; $i < 64; $i ++) {
//: my $b0 = $i * 8;
//: my $b1 = $i * 8 + 7;
//: &eperl::flop("-nodeclare  -norst -en \"dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[${i}]\" -d \"dat_out_bypass_data_w[${b1}:${b0}]\" -q dat_out_bypass_data[${b1}:${b0}]");
//: }
//:
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_pvld <= 1'b0;
   end else begin
       dat_out_pvld <= dat_out_pvld_w;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_flag <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld_w) == 1'b1) begin
           dat_out_flag <= dat_out_flag_w;
       // VCS coverage off
       end else if ((dat_out_pvld_w) == 1'b0) begin
       end else begin
           dat_out_flag <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dat_out_bypass_mask <= {64{1'b0}};
   end else begin
       if ((dat_out_bypass_p0_vld_w) == 1'b1) begin
           dat_out_bypass_mask <= dat_out_bypass_mask_w;
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w) == 1'b0) begin
       end else begin
           dat_out_bypass_mask <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[0]) == 1'b1) begin
           dat_out_bypass_data[7:0] <= dat_out_bypass_data_w[7:0];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[0]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[7:0] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[1]) == 1'b1) begin
           dat_out_bypass_data[15:8] <= dat_out_bypass_data_w[15:8];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[1]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[15:8] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[2]) == 1'b1) begin
           dat_out_bypass_data[23:16] <= dat_out_bypass_data_w[23:16];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[2]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[23:16] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[3]) == 1'b1) begin
           dat_out_bypass_data[31:24] <= dat_out_bypass_data_w[31:24];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[3]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[31:24] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[4]) == 1'b1) begin
           dat_out_bypass_data[39:32] <= dat_out_bypass_data_w[39:32];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[4]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[39:32] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[5]) == 1'b1) begin
           dat_out_bypass_data[47:40] <= dat_out_bypass_data_w[47:40];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[5]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[47:40] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[6]) == 1'b1) begin
           dat_out_bypass_data[55:48] <= dat_out_bypass_data_w[55:48];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[6]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[55:48] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[7]) == 1'b1) begin
           dat_out_bypass_data[63:56] <= dat_out_bypass_data_w[63:56];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[7]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[63:56] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[8]) == 1'b1) begin
           dat_out_bypass_data[71:64] <= dat_out_bypass_data_w[71:64];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[8]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[71:64] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[9]) == 1'b1) begin
           dat_out_bypass_data[79:72] <= dat_out_bypass_data_w[79:72];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[9]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[79:72] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[10]) == 1'b1) begin
           dat_out_bypass_data[87:80] <= dat_out_bypass_data_w[87:80];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[10]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[87:80] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[11]) == 1'b1) begin
           dat_out_bypass_data[95:88] <= dat_out_bypass_data_w[95:88];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[11]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[95:88] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[12]) == 1'b1) begin
           dat_out_bypass_data[103:96] <= dat_out_bypass_data_w[103:96];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[12]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[103:96] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[13]) == 1'b1) begin
           dat_out_bypass_data[111:104] <= dat_out_bypass_data_w[111:104];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[13]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[111:104] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[14]) == 1'b1) begin
           dat_out_bypass_data[119:112] <= dat_out_bypass_data_w[119:112];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[14]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[119:112] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[15]) == 1'b1) begin
           dat_out_bypass_data[127:120] <= dat_out_bypass_data_w[127:120];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[15]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[127:120] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[16]) == 1'b1) begin
           dat_out_bypass_data[135:128] <= dat_out_bypass_data_w[135:128];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[16]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[135:128] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[17]) == 1'b1) begin
           dat_out_bypass_data[143:136] <= dat_out_bypass_data_w[143:136];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[17]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[143:136] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[18]) == 1'b1) begin
           dat_out_bypass_data[151:144] <= dat_out_bypass_data_w[151:144];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[18]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[151:144] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[19]) == 1'b1) begin
           dat_out_bypass_data[159:152] <= dat_out_bypass_data_w[159:152];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[19]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[159:152] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[20]) == 1'b1) begin
           dat_out_bypass_data[167:160] <= dat_out_bypass_data_w[167:160];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[20]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[167:160] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[21]) == 1'b1) begin
           dat_out_bypass_data[175:168] <= dat_out_bypass_data_w[175:168];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[21]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[175:168] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[22]) == 1'b1) begin
           dat_out_bypass_data[183:176] <= dat_out_bypass_data_w[183:176];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[22]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[183:176] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[23]) == 1'b1) begin
           dat_out_bypass_data[191:184] <= dat_out_bypass_data_w[191:184];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[23]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[191:184] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[24]) == 1'b1) begin
           dat_out_bypass_data[199:192] <= dat_out_bypass_data_w[199:192];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[24]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[199:192] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[25]) == 1'b1) begin
           dat_out_bypass_data[207:200] <= dat_out_bypass_data_w[207:200];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[25]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[207:200] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[26]) == 1'b1) begin
           dat_out_bypass_data[215:208] <= dat_out_bypass_data_w[215:208];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[26]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[215:208] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[27]) == 1'b1) begin
           dat_out_bypass_data[223:216] <= dat_out_bypass_data_w[223:216];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[27]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[223:216] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[28]) == 1'b1) begin
           dat_out_bypass_data[231:224] <= dat_out_bypass_data_w[231:224];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[28]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[231:224] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[29]) == 1'b1) begin
           dat_out_bypass_data[239:232] <= dat_out_bypass_data_w[239:232];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[29]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[239:232] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[30]) == 1'b1) begin
           dat_out_bypass_data[247:240] <= dat_out_bypass_data_w[247:240];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[30]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[247:240] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[31]) == 1'b1) begin
           dat_out_bypass_data[255:248] <= dat_out_bypass_data_w[255:248];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[31]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[255:248] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[32]) == 1'b1) begin
           dat_out_bypass_data[263:256] <= dat_out_bypass_data_w[263:256];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[32]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[263:256] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[33]) == 1'b1) begin
           dat_out_bypass_data[271:264] <= dat_out_bypass_data_w[271:264];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[33]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[271:264] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[34]) == 1'b1) begin
           dat_out_bypass_data[279:272] <= dat_out_bypass_data_w[279:272];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[34]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[279:272] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[35]) == 1'b1) begin
           dat_out_bypass_data[287:280] <= dat_out_bypass_data_w[287:280];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[35]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[287:280] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[36]) == 1'b1) begin
           dat_out_bypass_data[295:288] <= dat_out_bypass_data_w[295:288];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[36]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[295:288] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[37]) == 1'b1) begin
           dat_out_bypass_data[303:296] <= dat_out_bypass_data_w[303:296];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[37]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[303:296] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[38]) == 1'b1) begin
           dat_out_bypass_data[311:304] <= dat_out_bypass_data_w[311:304];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[38]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[311:304] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[39]) == 1'b1) begin
           dat_out_bypass_data[319:312] <= dat_out_bypass_data_w[319:312];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[39]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[319:312] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[40]) == 1'b1) begin
           dat_out_bypass_data[327:320] <= dat_out_bypass_data_w[327:320];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[40]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[327:320] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[41]) == 1'b1) begin
           dat_out_bypass_data[335:328] <= dat_out_bypass_data_w[335:328];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[41]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[335:328] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[42]) == 1'b1) begin
           dat_out_bypass_data[343:336] <= dat_out_bypass_data_w[343:336];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[42]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[343:336] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[43]) == 1'b1) begin
           dat_out_bypass_data[351:344] <= dat_out_bypass_data_w[351:344];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[43]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[351:344] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[44]) == 1'b1) begin
           dat_out_bypass_data[359:352] <= dat_out_bypass_data_w[359:352];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[44]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[359:352] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[45]) == 1'b1) begin
           dat_out_bypass_data[367:360] <= dat_out_bypass_data_w[367:360];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[45]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[367:360] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[46]) == 1'b1) begin
           dat_out_bypass_data[375:368] <= dat_out_bypass_data_w[375:368];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[46]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[375:368] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[47]) == 1'b1) begin
           dat_out_bypass_data[383:376] <= dat_out_bypass_data_w[383:376];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[47]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[383:376] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[48]) == 1'b1) begin
           dat_out_bypass_data[391:384] <= dat_out_bypass_data_w[391:384];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[48]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[391:384] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[49]) == 1'b1) begin
           dat_out_bypass_data[399:392] <= dat_out_bypass_data_w[399:392];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[49]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[399:392] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[50]) == 1'b1) begin
           dat_out_bypass_data[407:400] <= dat_out_bypass_data_w[407:400];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[50]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[407:400] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[51]) == 1'b1) begin
           dat_out_bypass_data[415:408] <= dat_out_bypass_data_w[415:408];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[51]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[415:408] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[52]) == 1'b1) begin
           dat_out_bypass_data[423:416] <= dat_out_bypass_data_w[423:416];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[52]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[423:416] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[53]) == 1'b1) begin
           dat_out_bypass_data[431:424] <= dat_out_bypass_data_w[431:424];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[53]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[431:424] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[54]) == 1'b1) begin
           dat_out_bypass_data[439:432] <= dat_out_bypass_data_w[439:432];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[54]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[439:432] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[55]) == 1'b1) begin
           dat_out_bypass_data[447:440] <= dat_out_bypass_data_w[447:440];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[55]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[447:440] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[56]) == 1'b1) begin
           dat_out_bypass_data[455:448] <= dat_out_bypass_data_w[455:448];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[56]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[455:448] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[57]) == 1'b1) begin
           dat_out_bypass_data[463:456] <= dat_out_bypass_data_w[463:456];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[57]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[463:456] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[58]) == 1'b1) begin
           dat_out_bypass_data[471:464] <= dat_out_bypass_data_w[471:464];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[58]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[471:464] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[59]) == 1'b1) begin
           dat_out_bypass_data[479:472] <= dat_out_bypass_data_w[479:472];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[59]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[479:472] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[60]) == 1'b1) begin
           dat_out_bypass_data[487:480] <= dat_out_bypass_data_w[487:480];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[60]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[487:480] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[61]) == 1'b1) begin
           dat_out_bypass_data[495:488] <= dat_out_bypass_data_w[495:488];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[61]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[495:488] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[62]) == 1'b1) begin
           dat_out_bypass_data[503:496] <= dat_out_bypass_data_w[503:496];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[62]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[503:496] <= 'bx;
       // VCS coverage on
       end
end
always @(posedge nvdla_core_clk) begin
       if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[63]) == 1'b1) begin
           dat_out_bypass_data[511:504] <= dat_out_bypass_data_w[511:504];
       // VCS coverage off
       end else if ((dat_out_bypass_p0_vld_w & dat_out_bypass_mask_w[63]) == 1'b0) begin
       end else begin
           dat_out_bypass_data[511:504] <= 'bx;
       // VCS coverage on
       end
end

//| eperl: generated_end (DO NOT EDIT ABOVE)

assign dat_out_wg_data = {512{1'b0}};
assign dat_out_wg_mask = {64{1'b0}};
//////////////////////////////////////////////////////////////
///// finial registers                                   /////
//////////////////////////////////////////////////////////////
assign dat_out_data = is_winograd_d1[20] ? dat_out_wg_data : dat_out_bypass_data;
assign dat_out_mask = ~dat_out_pvld ? 'b0 : is_winograd_d1[21] ? dat_out_wg_mask : dat_out_bypass_mask;
//: my $kk=64;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dat_out_pvld\" -q dl_out_pvld");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dat_out_pvld | dl_out_pvld\" -d \"dat_out_mask\" -q dl_out_mask");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dat_out_pvld\" -d \"dat_out_flag\" -q dl_out_flag");
//: my $i;
//: my $b0;
//: my $b1;
//: my $kk= 8;
//: for($i = 0; $i < 64; $i ++) {
//: $b0 = $i * 8;
//: $b1 = $i * 8 + 7;
//: &eperl::flop("-wid ${kk}  -norst -en \"dat_out_mask[$i]\" -d \"dat_out_data[${b1}:${b0}]\" -q dl_out_data${i}");
//: }
//: print "\n\n\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_pvld <= 1'b0;
   end else begin
       dl_out_pvld <= dat_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_mask <= {64{1'b0}};
   end else begin
       if ((dat_out_pvld | dl_out_pvld) == 1'b1) begin
           dl_out_mask <= dat_out_mask;
       // VCS coverage off
       end else if ((dat_out_pvld | dl_out_pvld) == 1'b0) begin
       end else begin
           dl_out_mask <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_flag <= {9{1'b0}};
   end else begin
       if ((dat_out_pvld) == 1'b1) begin
           dl_out_flag <= dat_out_flag;
       // VCS coverage off
       end else if ((dat_out_pvld) == 1'b0) begin
       end else begin
           dl_out_flag <= 'bx;
       // VCS coverage on
       end
   end
end
reg [7:0] dl_out_data0;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[0]) == 1'b1) begin
           dl_out_data0 <= dat_out_data[7:0];
       // VCS coverage off
       end else if ((dat_out_mask[0]) == 1'b0) begin
       end else begin
           dl_out_data0 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data1;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[1]) == 1'b1) begin
           dl_out_data1 <= dat_out_data[15:8];
       // VCS coverage off
       end else if ((dat_out_mask[1]) == 1'b0) begin
       end else begin
           dl_out_data1 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data2;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[2]) == 1'b1) begin
           dl_out_data2 <= dat_out_data[23:16];
       // VCS coverage off
       end else if ((dat_out_mask[2]) == 1'b0) begin
       end else begin
           dl_out_data2 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data3;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[3]) == 1'b1) begin
           dl_out_data3 <= dat_out_data[31:24];
       // VCS coverage off
       end else if ((dat_out_mask[3]) == 1'b0) begin
       end else begin
           dl_out_data3 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data4;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[4]) == 1'b1) begin
           dl_out_data4 <= dat_out_data[39:32];
       // VCS coverage off
       end else if ((dat_out_mask[4]) == 1'b0) begin
       end else begin
           dl_out_data4 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data5;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[5]) == 1'b1) begin
           dl_out_data5 <= dat_out_data[47:40];
       // VCS coverage off
       end else if ((dat_out_mask[5]) == 1'b0) begin
       end else begin
           dl_out_data5 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data6;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[6]) == 1'b1) begin
           dl_out_data6 <= dat_out_data[55:48];
       // VCS coverage off
       end else if ((dat_out_mask[6]) == 1'b0) begin
       end else begin
           dl_out_data6 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data7;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[7]) == 1'b1) begin
           dl_out_data7 <= dat_out_data[63:56];
       // VCS coverage off
       end else if ((dat_out_mask[7]) == 1'b0) begin
       end else begin
           dl_out_data7 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data8;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[8]) == 1'b1) begin
           dl_out_data8 <= dat_out_data[71:64];
       // VCS coverage off
       end else if ((dat_out_mask[8]) == 1'b0) begin
       end else begin
           dl_out_data8 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data9;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[9]) == 1'b1) begin
           dl_out_data9 <= dat_out_data[79:72];
       // VCS coverage off
       end else if ((dat_out_mask[9]) == 1'b0) begin
       end else begin
           dl_out_data9 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data10;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[10]) == 1'b1) begin
           dl_out_data10 <= dat_out_data[87:80];
       // VCS coverage off
       end else if ((dat_out_mask[10]) == 1'b0) begin
       end else begin
           dl_out_data10 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data11;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[11]) == 1'b1) begin
           dl_out_data11 <= dat_out_data[95:88];
       // VCS coverage off
       end else if ((dat_out_mask[11]) == 1'b0) begin
       end else begin
           dl_out_data11 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data12;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[12]) == 1'b1) begin
           dl_out_data12 <= dat_out_data[103:96];
       // VCS coverage off
       end else if ((dat_out_mask[12]) == 1'b0) begin
       end else begin
           dl_out_data12 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data13;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[13]) == 1'b1) begin
           dl_out_data13 <= dat_out_data[111:104];
       // VCS coverage off
       end else if ((dat_out_mask[13]) == 1'b0) begin
       end else begin
           dl_out_data13 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data14;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[14]) == 1'b1) begin
           dl_out_data14 <= dat_out_data[119:112];
       // VCS coverage off
       end else if ((dat_out_mask[14]) == 1'b0) begin
       end else begin
           dl_out_data14 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data15;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[15]) == 1'b1) begin
           dl_out_data15 <= dat_out_data[127:120];
       // VCS coverage off
       end else if ((dat_out_mask[15]) == 1'b0) begin
       end else begin
           dl_out_data15 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data16;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[16]) == 1'b1) begin
           dl_out_data16 <= dat_out_data[135:128];
       // VCS coverage off
       end else if ((dat_out_mask[16]) == 1'b0) begin
       end else begin
           dl_out_data16 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data17;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[17]) == 1'b1) begin
           dl_out_data17 <= dat_out_data[143:136];
       // VCS coverage off
       end else if ((dat_out_mask[17]) == 1'b0) begin
       end else begin
           dl_out_data17 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data18;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[18]) == 1'b1) begin
           dl_out_data18 <= dat_out_data[151:144];
       // VCS coverage off
       end else if ((dat_out_mask[18]) == 1'b0) begin
       end else begin
           dl_out_data18 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data19;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[19]) == 1'b1) begin
           dl_out_data19 <= dat_out_data[159:152];
       // VCS coverage off
       end else if ((dat_out_mask[19]) == 1'b0) begin
       end else begin
           dl_out_data19 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data20;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[20]) == 1'b1) begin
           dl_out_data20 <= dat_out_data[167:160];
       // VCS coverage off
       end else if ((dat_out_mask[20]) == 1'b0) begin
       end else begin
           dl_out_data20 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data21;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[21]) == 1'b1) begin
           dl_out_data21 <= dat_out_data[175:168];
       // VCS coverage off
       end else if ((dat_out_mask[21]) == 1'b0) begin
       end else begin
           dl_out_data21 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data22;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[22]) == 1'b1) begin
           dl_out_data22 <= dat_out_data[183:176];
       // VCS coverage off
       end else if ((dat_out_mask[22]) == 1'b0) begin
       end else begin
           dl_out_data22 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data23;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[23]) == 1'b1) begin
           dl_out_data23 <= dat_out_data[191:184];
       // VCS coverage off
       end else if ((dat_out_mask[23]) == 1'b0) begin
       end else begin
           dl_out_data23 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data24;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[24]) == 1'b1) begin
           dl_out_data24 <= dat_out_data[199:192];
       // VCS coverage off
       end else if ((dat_out_mask[24]) == 1'b0) begin
       end else begin
           dl_out_data24 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data25;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[25]) == 1'b1) begin
           dl_out_data25 <= dat_out_data[207:200];
       // VCS coverage off
       end else if ((dat_out_mask[25]) == 1'b0) begin
       end else begin
           dl_out_data25 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data26;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[26]) == 1'b1) begin
           dl_out_data26 <= dat_out_data[215:208];
       // VCS coverage off
       end else if ((dat_out_mask[26]) == 1'b0) begin
       end else begin
           dl_out_data26 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data27;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[27]) == 1'b1) begin
           dl_out_data27 <= dat_out_data[223:216];
       // VCS coverage off
       end else if ((dat_out_mask[27]) == 1'b0) begin
       end else begin
           dl_out_data27 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data28;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[28]) == 1'b1) begin
           dl_out_data28 <= dat_out_data[231:224];
       // VCS coverage off
       end else if ((dat_out_mask[28]) == 1'b0) begin
       end else begin
           dl_out_data28 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data29;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[29]) == 1'b1) begin
           dl_out_data29 <= dat_out_data[239:232];
       // VCS coverage off
       end else if ((dat_out_mask[29]) == 1'b0) begin
       end else begin
           dl_out_data29 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data30;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[30]) == 1'b1) begin
           dl_out_data30 <= dat_out_data[247:240];
       // VCS coverage off
       end else if ((dat_out_mask[30]) == 1'b0) begin
       end else begin
           dl_out_data30 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data31;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[31]) == 1'b1) begin
           dl_out_data31 <= dat_out_data[255:248];
       // VCS coverage off
       end else if ((dat_out_mask[31]) == 1'b0) begin
       end else begin
           dl_out_data31 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data32;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[32]) == 1'b1) begin
           dl_out_data32 <= dat_out_data[263:256];
       // VCS coverage off
       end else if ((dat_out_mask[32]) == 1'b0) begin
       end else begin
           dl_out_data32 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data33;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[33]) == 1'b1) begin
           dl_out_data33 <= dat_out_data[271:264];
       // VCS coverage off
       end else if ((dat_out_mask[33]) == 1'b0) begin
       end else begin
           dl_out_data33 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data34;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[34]) == 1'b1) begin
           dl_out_data34 <= dat_out_data[279:272];
       // VCS coverage off
       end else if ((dat_out_mask[34]) == 1'b0) begin
       end else begin
           dl_out_data34 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data35;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[35]) == 1'b1) begin
           dl_out_data35 <= dat_out_data[287:280];
       // VCS coverage off
       end else if ((dat_out_mask[35]) == 1'b0) begin
       end else begin
           dl_out_data35 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data36;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[36]) == 1'b1) begin
           dl_out_data36 <= dat_out_data[295:288];
       // VCS coverage off
       end else if ((dat_out_mask[36]) == 1'b0) begin
       end else begin
           dl_out_data36 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data37;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[37]) == 1'b1) begin
           dl_out_data37 <= dat_out_data[303:296];
       // VCS coverage off
       end else if ((dat_out_mask[37]) == 1'b0) begin
       end else begin
           dl_out_data37 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data38;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[38]) == 1'b1) begin
           dl_out_data38 <= dat_out_data[311:304];
       // VCS coverage off
       end else if ((dat_out_mask[38]) == 1'b0) begin
       end else begin
           dl_out_data38 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data39;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[39]) == 1'b1) begin
           dl_out_data39 <= dat_out_data[319:312];
       // VCS coverage off
       end else if ((dat_out_mask[39]) == 1'b0) begin
       end else begin
           dl_out_data39 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data40;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[40]) == 1'b1) begin
           dl_out_data40 <= dat_out_data[327:320];
       // VCS coverage off
       end else if ((dat_out_mask[40]) == 1'b0) begin
       end else begin
           dl_out_data40 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data41;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[41]) == 1'b1) begin
           dl_out_data41 <= dat_out_data[335:328];
       // VCS coverage off
       end else if ((dat_out_mask[41]) == 1'b0) begin
       end else begin
           dl_out_data41 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data42;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[42]) == 1'b1) begin
           dl_out_data42 <= dat_out_data[343:336];
       // VCS coverage off
       end else if ((dat_out_mask[42]) == 1'b0) begin
       end else begin
           dl_out_data42 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data43;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[43]) == 1'b1) begin
           dl_out_data43 <= dat_out_data[351:344];
       // VCS coverage off
       end else if ((dat_out_mask[43]) == 1'b0) begin
       end else begin
           dl_out_data43 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data44;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[44]) == 1'b1) begin
           dl_out_data44 <= dat_out_data[359:352];
       // VCS coverage off
       end else if ((dat_out_mask[44]) == 1'b0) begin
       end else begin
           dl_out_data44 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data45;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[45]) == 1'b1) begin
           dl_out_data45 <= dat_out_data[367:360];
       // VCS coverage off
       end else if ((dat_out_mask[45]) == 1'b0) begin
       end else begin
           dl_out_data45 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data46;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[46]) == 1'b1) begin
           dl_out_data46 <= dat_out_data[375:368];
       // VCS coverage off
       end else if ((dat_out_mask[46]) == 1'b0) begin
       end else begin
           dl_out_data46 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data47;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[47]) == 1'b1) begin
           dl_out_data47 <= dat_out_data[383:376];
       // VCS coverage off
       end else if ((dat_out_mask[47]) == 1'b0) begin
       end else begin
           dl_out_data47 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data48;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[48]) == 1'b1) begin
           dl_out_data48 <= dat_out_data[391:384];
       // VCS coverage off
       end else if ((dat_out_mask[48]) == 1'b0) begin
       end else begin
           dl_out_data48 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data49;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[49]) == 1'b1) begin
           dl_out_data49 <= dat_out_data[399:392];
       // VCS coverage off
       end else if ((dat_out_mask[49]) == 1'b0) begin
       end else begin
           dl_out_data49 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data50;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[50]) == 1'b1) begin
           dl_out_data50 <= dat_out_data[407:400];
       // VCS coverage off
       end else if ((dat_out_mask[50]) == 1'b0) begin
       end else begin
           dl_out_data50 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data51;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[51]) == 1'b1) begin
           dl_out_data51 <= dat_out_data[415:408];
       // VCS coverage off
       end else if ((dat_out_mask[51]) == 1'b0) begin
       end else begin
           dl_out_data51 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data52;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[52]) == 1'b1) begin
           dl_out_data52 <= dat_out_data[423:416];
       // VCS coverage off
       end else if ((dat_out_mask[52]) == 1'b0) begin
       end else begin
           dl_out_data52 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data53;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[53]) == 1'b1) begin
           dl_out_data53 <= dat_out_data[431:424];
       // VCS coverage off
       end else if ((dat_out_mask[53]) == 1'b0) begin
       end else begin
           dl_out_data53 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data54;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[54]) == 1'b1) begin
           dl_out_data54 <= dat_out_data[439:432];
       // VCS coverage off
       end else if ((dat_out_mask[54]) == 1'b0) begin
       end else begin
           dl_out_data54 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data55;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[55]) == 1'b1) begin
           dl_out_data55 <= dat_out_data[447:440];
       // VCS coverage off
       end else if ((dat_out_mask[55]) == 1'b0) begin
       end else begin
           dl_out_data55 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data56;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[56]) == 1'b1) begin
           dl_out_data56 <= dat_out_data[455:448];
       // VCS coverage off
       end else if ((dat_out_mask[56]) == 1'b0) begin
       end else begin
           dl_out_data56 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data57;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[57]) == 1'b1) begin
           dl_out_data57 <= dat_out_data[463:456];
       // VCS coverage off
       end else if ((dat_out_mask[57]) == 1'b0) begin
       end else begin
           dl_out_data57 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data58;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[58]) == 1'b1) begin
           dl_out_data58 <= dat_out_data[471:464];
       // VCS coverage off
       end else if ((dat_out_mask[58]) == 1'b0) begin
       end else begin
           dl_out_data58 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data59;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[59]) == 1'b1) begin
           dl_out_data59 <= dat_out_data[479:472];
       // VCS coverage off
       end else if ((dat_out_mask[59]) == 1'b0) begin
       end else begin
           dl_out_data59 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data60;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[60]) == 1'b1) begin
           dl_out_data60 <= dat_out_data[487:480];
       // VCS coverage off
       end else if ((dat_out_mask[60]) == 1'b0) begin
       end else begin
           dl_out_data60 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data61;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[61]) == 1'b1) begin
           dl_out_data61 <= dat_out_data[495:488];
       // VCS coverage off
       end else if ((dat_out_mask[61]) == 1'b0) begin
       end else begin
           dl_out_data61 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data62;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[62]) == 1'b1) begin
           dl_out_data62 <= dat_out_data[503:496];
       // VCS coverage off
       end else if ((dat_out_mask[62]) == 1'b0) begin
       end else begin
           dl_out_data62 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] dl_out_data63;
always @(posedge nvdla_core_clk) begin
       if ((dat_out_mask[63]) == 1'b1) begin
           dl_out_data63 <= dat_out_data[511:504];
       // VCS coverage off
       end else if ((dat_out_mask[63]) == 1'b0) begin
       end else begin
           dl_out_data63 <= 'bx;
       // VCS coverage on
       end
end




//| eperl: generated_end (DO NOT EDIT ABOVE)
//////////////////////////////////////////////////////////////
///// registers for retiming                             /////
//////////////////////////////////////////////////////////////
assign sc2mac_dat_pd_w = ~dl_out_pvld ? 9'b0 : dl_out_flag;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dl_out_pvld\" -q dl_out_pvld_d1");
//: my $kk=64;
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dl_out_pvld\" -q sc2mac_dat_a_pvld");
//: &eperl::flop("-nodeclare   -rval \"1'b0\"   -d \"dl_out_pvld\" -q sc2mac_dat_b_pvld");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"sc2mac_dat_pd_w\" -q sc2mac_dat_a_pd");
//: &eperl::flop("-nodeclare   -rval \"{9{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"sc2mac_dat_pd_w\" -q sc2mac_dat_b_pd");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"dl_out_mask\" -q sc2mac_dat_a_mask");
//: &eperl::flop("-nodeclare   -rval \"{${kk}{1'b0}}\"  -en \"dl_out_pvld | dl_out_pvld_d1\" -d \"dl_out_mask\" -q sc2mac_dat_b_mask");
//: my $i;
//: for($i = 0; $i < 64; $i ++) {
//: &eperl::flop("-wid 8 -norst -en \"dl_out_mask[${i}]\" -d \"dl_out_data${i}\" -q sc2mac_dat_a_data${i}");
//: }
//: print "\n\n";
//:
//: for($i = 0; $i < 64; $i ++) {
//: &eperl::flop("-wid 8  -norst -en \"dl_out_mask[${i}]\" -d \"dl_out_data${i}\" -q sc2mac_dat_b_data${i}");
//: }
//: print "\n\n";
//| eperl: generated_beg (DO NOT EDIT BELOW)
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       dl_out_pvld_d1 <= 1'b0;
   end else begin
       dl_out_pvld_d1 <= dl_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_a_pvld <= 1'b0;
   end else begin
       sc2mac_dat_a_pvld <= dl_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_b_pvld <= 1'b0;
   end else begin
       sc2mac_dat_b_pvld <= dl_out_pvld;
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_a_pd <= {9{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_a_pd <= sc2mac_dat_pd_w;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_a_pd <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_b_pd <= {9{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_b_pd <= sc2mac_dat_pd_w;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_b_pd <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_a_mask <= {64{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_a_mask <= dl_out_mask;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_a_mask <= 'bx;
       // VCS coverage on
       end
   end
end
always @(posedge nvdla_core_clk) begin
   if (!nvdla_core_rstn) begin
       sc2mac_dat_b_mask <= {64{1'b0}};
   end else begin
       if ((dl_out_pvld | dl_out_pvld_d1) == 1'b1) begin
           sc2mac_dat_b_mask <= dl_out_mask;
       // VCS coverage off
       end else if ((dl_out_pvld | dl_out_pvld_d1) == 1'b0) begin
       end else begin
           sc2mac_dat_b_mask <= 'bx;
       // VCS coverage on
       end
   end
end
reg [7:0] sc2mac_dat_a_data0;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[0]) == 1'b1) begin
           sc2mac_dat_a_data0 <= dl_out_data0;
       // VCS coverage off
       end else if ((dl_out_mask[0]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data0 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data1;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[1]) == 1'b1) begin
           sc2mac_dat_a_data1 <= dl_out_data1;
       // VCS coverage off
       end else if ((dl_out_mask[1]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data1 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data2;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[2]) == 1'b1) begin
           sc2mac_dat_a_data2 <= dl_out_data2;
       // VCS coverage off
       end else if ((dl_out_mask[2]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data2 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data3;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[3]) == 1'b1) begin
           sc2mac_dat_a_data3 <= dl_out_data3;
       // VCS coverage off
       end else if ((dl_out_mask[3]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data3 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data4;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[4]) == 1'b1) begin
           sc2mac_dat_a_data4 <= dl_out_data4;
       // VCS coverage off
       end else if ((dl_out_mask[4]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data4 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data5;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[5]) == 1'b1) begin
           sc2mac_dat_a_data5 <= dl_out_data5;
       // VCS coverage off
       end else if ((dl_out_mask[5]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data5 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data6;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[6]) == 1'b1) begin
           sc2mac_dat_a_data6 <= dl_out_data6;
       // VCS coverage off
       end else if ((dl_out_mask[6]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data6 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data7;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[7]) == 1'b1) begin
           sc2mac_dat_a_data7 <= dl_out_data7;
       // VCS coverage off
       end else if ((dl_out_mask[7]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data7 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data8;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[8]) == 1'b1) begin
           sc2mac_dat_a_data8 <= dl_out_data8;
       // VCS coverage off
       end else if ((dl_out_mask[8]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data8 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data9;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[9]) == 1'b1) begin
           sc2mac_dat_a_data9 <= dl_out_data9;
       // VCS coverage off
       end else if ((dl_out_mask[9]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data9 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data10;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[10]) == 1'b1) begin
           sc2mac_dat_a_data10 <= dl_out_data10;
       // VCS coverage off
       end else if ((dl_out_mask[10]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data10 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data11;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[11]) == 1'b1) begin
           sc2mac_dat_a_data11 <= dl_out_data11;
       // VCS coverage off
       end else if ((dl_out_mask[11]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data11 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data12;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[12]) == 1'b1) begin
           sc2mac_dat_a_data12 <= dl_out_data12;
       // VCS coverage off
       end else if ((dl_out_mask[12]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data12 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data13;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[13]) == 1'b1) begin
           sc2mac_dat_a_data13 <= dl_out_data13;
       // VCS coverage off
       end else if ((dl_out_mask[13]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data13 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data14;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[14]) == 1'b1) begin
           sc2mac_dat_a_data14 <= dl_out_data14;
       // VCS coverage off
       end else if ((dl_out_mask[14]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data14 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data15;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[15]) == 1'b1) begin
           sc2mac_dat_a_data15 <= dl_out_data15;
       // VCS coverage off
       end else if ((dl_out_mask[15]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data15 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data16;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[16]) == 1'b1) begin
           sc2mac_dat_a_data16 <= dl_out_data16;
       // VCS coverage off
       end else if ((dl_out_mask[16]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data16 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data17;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[17]) == 1'b1) begin
           sc2mac_dat_a_data17 <= dl_out_data17;
       // VCS coverage off
       end else if ((dl_out_mask[17]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data17 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data18;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[18]) == 1'b1) begin
           sc2mac_dat_a_data18 <= dl_out_data18;
       // VCS coverage off
       end else if ((dl_out_mask[18]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data18 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data19;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[19]) == 1'b1) begin
           sc2mac_dat_a_data19 <= dl_out_data19;
       // VCS coverage off
       end else if ((dl_out_mask[19]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data19 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data20;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[20]) == 1'b1) begin
           sc2mac_dat_a_data20 <= dl_out_data20;
       // VCS coverage off
       end else if ((dl_out_mask[20]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data20 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data21;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[21]) == 1'b1) begin
           sc2mac_dat_a_data21 <= dl_out_data21;
       // VCS coverage off
       end else if ((dl_out_mask[21]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data21 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data22;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[22]) == 1'b1) begin
           sc2mac_dat_a_data22 <= dl_out_data22;
       // VCS coverage off
       end else if ((dl_out_mask[22]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data22 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data23;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[23]) == 1'b1) begin
           sc2mac_dat_a_data23 <= dl_out_data23;
       // VCS coverage off
       end else if ((dl_out_mask[23]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data23 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data24;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[24]) == 1'b1) begin
           sc2mac_dat_a_data24 <= dl_out_data24;
       // VCS coverage off
       end else if ((dl_out_mask[24]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data24 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data25;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[25]) == 1'b1) begin
           sc2mac_dat_a_data25 <= dl_out_data25;
       // VCS coverage off
       end else if ((dl_out_mask[25]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data25 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data26;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[26]) == 1'b1) begin
           sc2mac_dat_a_data26 <= dl_out_data26;
       // VCS coverage off
       end else if ((dl_out_mask[26]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data26 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data27;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[27]) == 1'b1) begin
           sc2mac_dat_a_data27 <= dl_out_data27;
       // VCS coverage off
       end else if ((dl_out_mask[27]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data27 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data28;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[28]) == 1'b1) begin
           sc2mac_dat_a_data28 <= dl_out_data28;
       // VCS coverage off
       end else if ((dl_out_mask[28]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data28 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data29;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[29]) == 1'b1) begin
           sc2mac_dat_a_data29 <= dl_out_data29;
       // VCS coverage off
       end else if ((dl_out_mask[29]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data29 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data30;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[30]) == 1'b1) begin
           sc2mac_dat_a_data30 <= dl_out_data30;
       // VCS coverage off
       end else if ((dl_out_mask[30]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data30 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data31;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[31]) == 1'b1) begin
           sc2mac_dat_a_data31 <= dl_out_data31;
       // VCS coverage off
       end else if ((dl_out_mask[31]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data31 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data32;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[32]) == 1'b1) begin
           sc2mac_dat_a_data32 <= dl_out_data32;
       // VCS coverage off
       end else if ((dl_out_mask[32]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data32 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data33;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[33]) == 1'b1) begin
           sc2mac_dat_a_data33 <= dl_out_data33;
       // VCS coverage off
       end else if ((dl_out_mask[33]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data33 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data34;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[34]) == 1'b1) begin
           sc2mac_dat_a_data34 <= dl_out_data34;
       // VCS coverage off
       end else if ((dl_out_mask[34]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data34 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data35;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[35]) == 1'b1) begin
           sc2mac_dat_a_data35 <= dl_out_data35;
       // VCS coverage off
       end else if ((dl_out_mask[35]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data35 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data36;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[36]) == 1'b1) begin
           sc2mac_dat_a_data36 <= dl_out_data36;
       // VCS coverage off
       end else if ((dl_out_mask[36]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data36 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data37;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[37]) == 1'b1) begin
           sc2mac_dat_a_data37 <= dl_out_data37;
       // VCS coverage off
       end else if ((dl_out_mask[37]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data37 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data38;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[38]) == 1'b1) begin
           sc2mac_dat_a_data38 <= dl_out_data38;
       // VCS coverage off
       end else if ((dl_out_mask[38]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data38 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data39;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[39]) == 1'b1) begin
           sc2mac_dat_a_data39 <= dl_out_data39;
       // VCS coverage off
       end else if ((dl_out_mask[39]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data39 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data40;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[40]) == 1'b1) begin
           sc2mac_dat_a_data40 <= dl_out_data40;
       // VCS coverage off
       end else if ((dl_out_mask[40]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data40 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data41;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[41]) == 1'b1) begin
           sc2mac_dat_a_data41 <= dl_out_data41;
       // VCS coverage off
       end else if ((dl_out_mask[41]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data41 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data42;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[42]) == 1'b1) begin
           sc2mac_dat_a_data42 <= dl_out_data42;
       // VCS coverage off
       end else if ((dl_out_mask[42]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data42 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data43;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[43]) == 1'b1) begin
           sc2mac_dat_a_data43 <= dl_out_data43;
       // VCS coverage off
       end else if ((dl_out_mask[43]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data43 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data44;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[44]) == 1'b1) begin
           sc2mac_dat_a_data44 <= dl_out_data44;
       // VCS coverage off
       end else if ((dl_out_mask[44]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data44 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data45;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[45]) == 1'b1) begin
           sc2mac_dat_a_data45 <= dl_out_data45;
       // VCS coverage off
       end else if ((dl_out_mask[45]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data45 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data46;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[46]) == 1'b1) begin
           sc2mac_dat_a_data46 <= dl_out_data46;
       // VCS coverage off
       end else if ((dl_out_mask[46]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data46 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data47;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[47]) == 1'b1) begin
           sc2mac_dat_a_data47 <= dl_out_data47;
       // VCS coverage off
       end else if ((dl_out_mask[47]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data47 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data48;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[48]) == 1'b1) begin
           sc2mac_dat_a_data48 <= dl_out_data48;
       // VCS coverage off
       end else if ((dl_out_mask[48]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data48 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data49;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[49]) == 1'b1) begin
           sc2mac_dat_a_data49 <= dl_out_data49;
       // VCS coverage off
       end else if ((dl_out_mask[49]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data49 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data50;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[50]) == 1'b1) begin
           sc2mac_dat_a_data50 <= dl_out_data50;
       // VCS coverage off
       end else if ((dl_out_mask[50]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data50 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data51;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[51]) == 1'b1) begin
           sc2mac_dat_a_data51 <= dl_out_data51;
       // VCS coverage off
       end else if ((dl_out_mask[51]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data51 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data52;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[52]) == 1'b1) begin
           sc2mac_dat_a_data52 <= dl_out_data52;
       // VCS coverage off
       end else if ((dl_out_mask[52]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data52 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data53;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[53]) == 1'b1) begin
           sc2mac_dat_a_data53 <= dl_out_data53;
       // VCS coverage off
       end else if ((dl_out_mask[53]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data53 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data54;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[54]) == 1'b1) begin
           sc2mac_dat_a_data54 <= dl_out_data54;
       // VCS coverage off
       end else if ((dl_out_mask[54]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data54 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data55;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[55]) == 1'b1) begin
           sc2mac_dat_a_data55 <= dl_out_data55;
       // VCS coverage off
       end else if ((dl_out_mask[55]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data55 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data56;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[56]) == 1'b1) begin
           sc2mac_dat_a_data56 <= dl_out_data56;
       // VCS coverage off
       end else if ((dl_out_mask[56]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data56 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data57;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[57]) == 1'b1) begin
           sc2mac_dat_a_data57 <= dl_out_data57;
       // VCS coverage off
       end else if ((dl_out_mask[57]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data57 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data58;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[58]) == 1'b1) begin
           sc2mac_dat_a_data58 <= dl_out_data58;
       // VCS coverage off
       end else if ((dl_out_mask[58]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data58 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data59;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[59]) == 1'b1) begin
           sc2mac_dat_a_data59 <= dl_out_data59;
       // VCS coverage off
       end else if ((dl_out_mask[59]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data59 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data60;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[60]) == 1'b1) begin
           sc2mac_dat_a_data60 <= dl_out_data60;
       // VCS coverage off
       end else if ((dl_out_mask[60]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data60 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data61;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[61]) == 1'b1) begin
           sc2mac_dat_a_data61 <= dl_out_data61;
       // VCS coverage off
       end else if ((dl_out_mask[61]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data61 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data62;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[62]) == 1'b1) begin
           sc2mac_dat_a_data62 <= dl_out_data62;
       // VCS coverage off
       end else if ((dl_out_mask[62]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data62 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_a_data63;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[63]) == 1'b1) begin
           sc2mac_dat_a_data63 <= dl_out_data63;
       // VCS coverage off
       end else if ((dl_out_mask[63]) == 1'b0) begin
       end else begin
           sc2mac_dat_a_data63 <= 'bx;
       // VCS coverage on
       end
end


reg [7:0] sc2mac_dat_b_data0;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[0]) == 1'b1) begin
           sc2mac_dat_b_data0 <= dl_out_data0;
       // VCS coverage off
       end else if ((dl_out_mask[0]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data0 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data1;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[1]) == 1'b1) begin
           sc2mac_dat_b_data1 <= dl_out_data1;
       // VCS coverage off
       end else if ((dl_out_mask[1]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data1 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data2;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[2]) == 1'b1) begin
           sc2mac_dat_b_data2 <= dl_out_data2;
       // VCS coverage off
       end else if ((dl_out_mask[2]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data2 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data3;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[3]) == 1'b1) begin
           sc2mac_dat_b_data3 <= dl_out_data3;
       // VCS coverage off
       end else if ((dl_out_mask[3]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data3 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data4;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[4]) == 1'b1) begin
           sc2mac_dat_b_data4 <= dl_out_data4;
       // VCS coverage off
       end else if ((dl_out_mask[4]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data4 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data5;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[5]) == 1'b1) begin
           sc2mac_dat_b_data5 <= dl_out_data5;
       // VCS coverage off
       end else if ((dl_out_mask[5]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data5 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data6;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[6]) == 1'b1) begin
           sc2mac_dat_b_data6 <= dl_out_data6;
       // VCS coverage off
       end else if ((dl_out_mask[6]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data6 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data7;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[7]) == 1'b1) begin
           sc2mac_dat_b_data7 <= dl_out_data7;
       // VCS coverage off
       end else if ((dl_out_mask[7]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data7 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data8;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[8]) == 1'b1) begin
           sc2mac_dat_b_data8 <= dl_out_data8;
       // VCS coverage off
       end else if ((dl_out_mask[8]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data8 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data9;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[9]) == 1'b1) begin
           sc2mac_dat_b_data9 <= dl_out_data9;
       // VCS coverage off
       end else if ((dl_out_mask[9]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data9 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data10;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[10]) == 1'b1) begin
           sc2mac_dat_b_data10 <= dl_out_data10;
       // VCS coverage off
       end else if ((dl_out_mask[10]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data10 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data11;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[11]) == 1'b1) begin
           sc2mac_dat_b_data11 <= dl_out_data11;
       // VCS coverage off
       end else if ((dl_out_mask[11]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data11 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data12;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[12]) == 1'b1) begin
           sc2mac_dat_b_data12 <= dl_out_data12;
       // VCS coverage off
       end else if ((dl_out_mask[12]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data12 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data13;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[13]) == 1'b1) begin
           sc2mac_dat_b_data13 <= dl_out_data13;
       // VCS coverage off
       end else if ((dl_out_mask[13]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data13 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data14;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[14]) == 1'b1) begin
           sc2mac_dat_b_data14 <= dl_out_data14;
       // VCS coverage off
       end else if ((dl_out_mask[14]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data14 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data15;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[15]) == 1'b1) begin
           sc2mac_dat_b_data15 <= dl_out_data15;
       // VCS coverage off
       end else if ((dl_out_mask[15]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data15 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data16;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[16]) == 1'b1) begin
           sc2mac_dat_b_data16 <= dl_out_data16;
       // VCS coverage off
       end else if ((dl_out_mask[16]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data16 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data17;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[17]) == 1'b1) begin
           sc2mac_dat_b_data17 <= dl_out_data17;
       // VCS coverage off
       end else if ((dl_out_mask[17]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data17 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data18;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[18]) == 1'b1) begin
           sc2mac_dat_b_data18 <= dl_out_data18;
       // VCS coverage off
       end else if ((dl_out_mask[18]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data18 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data19;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[19]) == 1'b1) begin
           sc2mac_dat_b_data19 <= dl_out_data19;
       // VCS coverage off
       end else if ((dl_out_mask[19]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data19 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data20;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[20]) == 1'b1) begin
           sc2mac_dat_b_data20 <= dl_out_data20;
       // VCS coverage off
       end else if ((dl_out_mask[20]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data20 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data21;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[21]) == 1'b1) begin
           sc2mac_dat_b_data21 <= dl_out_data21;
       // VCS coverage off
       end else if ((dl_out_mask[21]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data21 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data22;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[22]) == 1'b1) begin
           sc2mac_dat_b_data22 <= dl_out_data22;
       // VCS coverage off
       end else if ((dl_out_mask[22]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data22 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data23;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[23]) == 1'b1) begin
           sc2mac_dat_b_data23 <= dl_out_data23;
       // VCS coverage off
       end else if ((dl_out_mask[23]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data23 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data24;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[24]) == 1'b1) begin
           sc2mac_dat_b_data24 <= dl_out_data24;
       // VCS coverage off
       end else if ((dl_out_mask[24]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data24 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data25;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[25]) == 1'b1) begin
           sc2mac_dat_b_data25 <= dl_out_data25;
       // VCS coverage off
       end else if ((dl_out_mask[25]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data25 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data26;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[26]) == 1'b1) begin
           sc2mac_dat_b_data26 <= dl_out_data26;
       // VCS coverage off
       end else if ((dl_out_mask[26]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data26 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data27;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[27]) == 1'b1) begin
           sc2mac_dat_b_data27 <= dl_out_data27;
       // VCS coverage off
       end else if ((dl_out_mask[27]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data27 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data28;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[28]) == 1'b1) begin
           sc2mac_dat_b_data28 <= dl_out_data28;
       // VCS coverage off
       end else if ((dl_out_mask[28]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data28 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data29;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[29]) == 1'b1) begin
           sc2mac_dat_b_data29 <= dl_out_data29;
       // VCS coverage off
       end else if ((dl_out_mask[29]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data29 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data30;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[30]) == 1'b1) begin
           sc2mac_dat_b_data30 <= dl_out_data30;
       // VCS coverage off
       end else if ((dl_out_mask[30]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data30 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data31;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[31]) == 1'b1) begin
           sc2mac_dat_b_data31 <= dl_out_data31;
       // VCS coverage off
       end else if ((dl_out_mask[31]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data31 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data32;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[32]) == 1'b1) begin
           sc2mac_dat_b_data32 <= dl_out_data32;
       // VCS coverage off
       end else if ((dl_out_mask[32]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data32 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data33;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[33]) == 1'b1) begin
           sc2mac_dat_b_data33 <= dl_out_data33;
       // VCS coverage off
       end else if ((dl_out_mask[33]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data33 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data34;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[34]) == 1'b1) begin
           sc2mac_dat_b_data34 <= dl_out_data34;
       // VCS coverage off
       end else if ((dl_out_mask[34]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data34 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data35;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[35]) == 1'b1) begin
           sc2mac_dat_b_data35 <= dl_out_data35;
       // VCS coverage off
       end else if ((dl_out_mask[35]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data35 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data36;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[36]) == 1'b1) begin
           sc2mac_dat_b_data36 <= dl_out_data36;
       // VCS coverage off
       end else if ((dl_out_mask[36]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data36 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data37;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[37]) == 1'b1) begin
           sc2mac_dat_b_data37 <= dl_out_data37;
       // VCS coverage off
       end else if ((dl_out_mask[37]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data37 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data38;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[38]) == 1'b1) begin
           sc2mac_dat_b_data38 <= dl_out_data38;
       // VCS coverage off
       end else if ((dl_out_mask[38]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data38 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data39;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[39]) == 1'b1) begin
           sc2mac_dat_b_data39 <= dl_out_data39;
       // VCS coverage off
       end else if ((dl_out_mask[39]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data39 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data40;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[40]) == 1'b1) begin
           sc2mac_dat_b_data40 <= dl_out_data40;
       // VCS coverage off
       end else if ((dl_out_mask[40]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data40 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data41;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[41]) == 1'b1) begin
           sc2mac_dat_b_data41 <= dl_out_data41;
       // VCS coverage off
       end else if ((dl_out_mask[41]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data41 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data42;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[42]) == 1'b1) begin
           sc2mac_dat_b_data42 <= dl_out_data42;
       // VCS coverage off
       end else if ((dl_out_mask[42]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data42 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data43;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[43]) == 1'b1) begin
           sc2mac_dat_b_data43 <= dl_out_data43;
       // VCS coverage off
       end else if ((dl_out_mask[43]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data43 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data44;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[44]) == 1'b1) begin
           sc2mac_dat_b_data44 <= dl_out_data44;
       // VCS coverage off
       end else if ((dl_out_mask[44]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data44 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data45;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[45]) == 1'b1) begin
           sc2mac_dat_b_data45 <= dl_out_data45;
       // VCS coverage off
       end else if ((dl_out_mask[45]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data45 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data46;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[46]) == 1'b1) begin
           sc2mac_dat_b_data46 <= dl_out_data46;
       // VCS coverage off
       end else if ((dl_out_mask[46]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data46 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data47;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[47]) == 1'b1) begin
           sc2mac_dat_b_data47 <= dl_out_data47;
       // VCS coverage off
       end else if ((dl_out_mask[47]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data47 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data48;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[48]) == 1'b1) begin
           sc2mac_dat_b_data48 <= dl_out_data48;
       // VCS coverage off
       end else if ((dl_out_mask[48]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data48 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data49;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[49]) == 1'b1) begin
           sc2mac_dat_b_data49 <= dl_out_data49;
       // VCS coverage off
       end else if ((dl_out_mask[49]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data49 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data50;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[50]) == 1'b1) begin
           sc2mac_dat_b_data50 <= dl_out_data50;
       // VCS coverage off
       end else if ((dl_out_mask[50]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data50 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data51;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[51]) == 1'b1) begin
           sc2mac_dat_b_data51 <= dl_out_data51;
       // VCS coverage off
       end else if ((dl_out_mask[51]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data51 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data52;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[52]) == 1'b1) begin
           sc2mac_dat_b_data52 <= dl_out_data52;
       // VCS coverage off
       end else if ((dl_out_mask[52]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data52 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data53;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[53]) == 1'b1) begin
           sc2mac_dat_b_data53 <= dl_out_data53;
       // VCS coverage off
       end else if ((dl_out_mask[53]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data53 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data54;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[54]) == 1'b1) begin
           sc2mac_dat_b_data54 <= dl_out_data54;
       // VCS coverage off
       end else if ((dl_out_mask[54]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data54 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data55;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[55]) == 1'b1) begin
           sc2mac_dat_b_data55 <= dl_out_data55;
       // VCS coverage off
       end else if ((dl_out_mask[55]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data55 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data56;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[56]) == 1'b1) begin
           sc2mac_dat_b_data56 <= dl_out_data56;
       // VCS coverage off
       end else if ((dl_out_mask[56]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data56 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data57;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[57]) == 1'b1) begin
           sc2mac_dat_b_data57 <= dl_out_data57;
       // VCS coverage off
       end else if ((dl_out_mask[57]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data57 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data58;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[58]) == 1'b1) begin
           sc2mac_dat_b_data58 <= dl_out_data58;
       // VCS coverage off
       end else if ((dl_out_mask[58]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data58 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data59;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[59]) == 1'b1) begin
           sc2mac_dat_b_data59 <= dl_out_data59;
       // VCS coverage off
       end else if ((dl_out_mask[59]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data59 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data60;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[60]) == 1'b1) begin
           sc2mac_dat_b_data60 <= dl_out_data60;
       // VCS coverage off
       end else if ((dl_out_mask[60]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data60 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data61;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[61]) == 1'b1) begin
           sc2mac_dat_b_data61 <= dl_out_data61;
       // VCS coverage off
       end else if ((dl_out_mask[61]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data61 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data62;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[62]) == 1'b1) begin
           sc2mac_dat_b_data62 <= dl_out_data62;
       // VCS coverage off
       end else if ((dl_out_mask[62]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data62 <= 'bx;
       // VCS coverage on
       end
end
reg [7:0] sc2mac_dat_b_data63;
always @(posedge nvdla_core_clk) begin
       if ((dl_out_mask[63]) == 1'b1) begin
           sc2mac_dat_b_data63 <= dl_out_data63;
       // VCS coverage off
       end else if ((dl_out_mask[63]) == 1'b0) begin
       end else begin
           sc2mac_dat_b_data63 <= 'bx;
       // VCS coverage on
       end
end


endmodule // NV_NVDLA_CSC_dl

module NV_soDLA_CSC_dl_for_check( // @[:@3.2]
  input          clock, // @[:@4.4]
  input          reset, // @[:@5.4]
  input          io_nvdla_core_clk, // @[:@6.4]
  input          io_nvdla_core_ng_clk, // @[:@6.4]
  input          io_nvdla_core_rstn, // @[:@6.4]
  input  [1:0]   io_sc_state, // @[:@6.4]
  input          io_sg2dl_pd_valid, // @[:@6.4]
  input  [30:0]  io_sg2dl_pd_bits, // @[:@6.4]
  input          io_sg2dl_reuse_rls, // @[:@6.4]
  input          io_cdma2sc_dat_updt_valid, // @[:@6.4]
  input  [14:0]  io_cdma2sc_dat_updt_bits_entries, // @[:@6.4]
  input  [13:0]  io_cdma2sc_dat_updt_bits_slices, // @[:@6.4]
  input          io_sc2cdma_dat_pending_req, // @[:@6.4]
  output         io_sc2cdma_dat_updt_valid, // @[:@6.4]
  output [14:0]  io_sc2cdma_dat_updt_bits_entries, // @[:@6.4]
  output [13:0]  io_sc2cdma_dat_updt_bits_slices, // @[:@6.4]
  output         io_sc2buf_dat_rd_addr_valid, // @[:@6.4]
  output [12:0]  io_sc2buf_dat_rd_addr_bits, // @[:@6.4]
  input          io_sc2buf_dat_rd_data_valid, // @[:@6.4]
  input  [511:0] io_sc2buf_dat_rd_data_bits, // @[:@6.4]
  output         io_sc2mac_dat_a_pvld, // @[:@6.4]
  output [63:0]  io_sc2mac_dat_a_mask, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_0, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_1, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_2, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_3, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_4, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_5, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_6, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_7, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_8, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_9, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_10, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_11, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_12, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_13, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_14, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_15, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_16, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_17, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_18, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_19, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_20, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_21, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_22, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_23, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_24, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_25, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_26, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_27, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_28, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_29, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_30, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_31, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_32, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_33, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_34, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_35, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_36, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_37, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_38, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_39, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_40, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_41, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_42, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_43, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_44, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_45, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_46, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_47, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_48, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_49, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_50, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_51, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_52, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_53, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_54, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_55, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_56, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_57, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_58, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_59, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_60, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_61, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_62, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_a_data_63, // @[:@6.4]
  output [8:0]   io_sc2mac_dat_a_pd, // @[:@6.4]
  output         io_sc2mac_dat_b_pvld, // @[:@6.4]
  output [63:0]  io_sc2mac_dat_b_mask, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_0, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_1, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_2, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_3, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_4, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_5, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_6, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_7, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_8, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_9, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_10, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_11, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_12, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_13, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_14, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_15, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_16, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_17, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_18, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_19, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_20, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_21, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_22, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_23, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_24, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_25, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_26, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_27, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_28, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_29, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_30, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_31, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_32, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_33, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_34, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_35, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_36, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_37, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_38, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_39, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_40, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_41, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_42, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_43, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_44, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_45, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_46, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_47, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_48, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_49, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_50, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_51, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_52, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_53, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_54, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_55, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_56, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_57, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_58, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_59, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_60, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_61, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_62, // @[:@6.4]
  output [7:0]   io_sc2mac_dat_b_data_63, // @[:@6.4]
  output [8:0]   io_sc2mac_dat_b_pd, // @[:@6.4]
  input          io_reg2dp_op_en, // @[:@6.4]
  input          io_reg2dp_conv_mode, // @[:@6.4]
  input  [4:0]   io_reg2dp_batches, // @[:@6.4]
  input  [1:0]   io_reg2dp_proc_precision, // @[:@6.4]
  input          io_reg2dp_datain_format, // @[:@6.4]
  input          io_reg2dp_skip_data_rls, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_channel_ext, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_height_ext, // @[:@6.4]
  input  [12:0]  io_reg2dp_datain_width_ext, // @[:@6.4]
  input  [1:0]   io_reg2dp_y_extension, // @[:@6.4]
  input  [12:0]  io_reg2dp_weight_channel_ext, // @[:@6.4]
  input  [13:0]  io_reg2dp_entries, // @[:@6.4]
  input  [12:0]  io_reg2dp_dataout_width, // @[:@6.4]
  input  [11:0]  io_reg2dp_rls_slices, // @[:@6.4]
  input  [2:0]   io_reg2dp_conv_x_stride_ext, // @[:@6.4]
  input  [2:0]   io_reg2dp_conv_y_stride_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_x_dilation_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_y_dilation_ext, // @[:@6.4]
  input  [4:0]   io_reg2dp_pad_left, // @[:@6.4]
  input  [4:0]   io_reg2dp_pad_top, // @[:@6.4]
  input  [15:0]  io_reg2dp_pad_value, // @[:@6.4]
  input  [4:0]   io_reg2dp_data_bank, // @[:@6.4]
  input  [1:0]   io_reg2dp_pra_truncate, // @[:@6.4]
  output         io_slcg_wg_en // @[:@6.4]
);
  wire  _T_207; // @[NV_NVDLA_CSC_dl_for_check.scala 81:38:@8.4]
  wire  is_sg_idle; // @[NV_NVDLA_CSC_dl_for_check.scala 85:31:@9.4]
  wire  is_sg_done; // @[NV_NVDLA_CSC_dl_for_check.scala 87:31:@11.4]
  wire  layer_st; // @[NV_NVDLA_CSC_dl_for_check.scala 94:32:@14.4]
  wire  is_conv; // @[NV_NVDLA_CSC_dl_for_check.scala 96:35:@16.4]
  wire  is_img; // @[NV_NVDLA_CSC_dl_for_check.scala 97:22:@17.4]
  wire [6:0] _T_216; // @[NV_NVDLA_CSC_dl_for_check.scala 105:53:@18.4]
  wire [6:0] _T_218; // @[NV_NVDLA_CSC_dl_for_check.scala 105:24:@19.4]
  wire [2:0] sub_h_total_w; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@20.4]
  wire [2:0] sub_h_cmp_w; // @[NV_NVDLA_CSC_dl_for_check.scala 106:22:@21.4]
  wire [3:0] _T_221; // @[NV_NVDLA_CSC_dl_for_check.scala 107:34:@22.4]
  wire [3:0] dataout_w_init; // @[NV_NVDLA_CSC_dl_for_check.scala 107:34:@23.4]
  wire [3:0] conv_x_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 108:73:@24.4]
  wire [1:0] _T_225; // @[NV_NVDLA_CSC_dl_for_check.scala 109:62:@26.4]
  wire [5:0] _T_228; // @[Cat.scala 30:58:@27.4]
  wire [4:0] _T_231; // @[Cat.scala 30:58:@28.4]
  wire [4:0] _GEN_681; // @[NV_NVDLA_CSC_dl_for_check.scala 111:74:@29.4]
  wire [5:0] _T_232; // @[NV_NVDLA_CSC_dl_for_check.scala 111:74:@29.4]
  wire  _T_233; // @[Mux.scala 46:19:@30.4]
  wire [5:0] _T_234; // @[Mux.scala 46:16:@31.4]
  wire  _T_235; // @[Mux.scala 46:19:@32.4]
  wire [5:0] pixel_x_stride_w; // @[Mux.scala 46:16:@33.4]
  wire  _T_237; // @[NV_NVDLA_CSC_dl_for_check.scala 113:88:@34.4]
  wire [5:0] _T_243; // @[NV_NVDLA_CSC_dl_for_check.scala 113:172:@36.4]
  wire [5:0] _T_244; // @[NV_NVDLA_CSC_dl_for_check.scala 113:58:@37.4]
  wire [6:0] _T_247; // @[Cat.scala 30:58:@38.4]
  wire [6:0] _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 114:81:@39.4]
  wire [7:0] _T_248; // @[NV_NVDLA_CSC_dl_for_check.scala 114:81:@39.4]
  wire [6:0] _T_249; // @[NV_NVDLA_CSC_dl_for_check.scala 114:81:@40.4]
  wire [6:0] _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 114:100:@42.4]
  wire [7:0] _T_251; // @[NV_NVDLA_CSC_dl_for_check.scala 114:100:@42.4]
  wire [6:0] _T_252; // @[NV_NVDLA_CSC_dl_for_check.scala 114:100:@43.4]
  wire [6:0] _T_255; // @[NV_NVDLA_CSC_dl_for_check.scala 115:58:@45.4]
  wire [5:0] _T_256; // @[NV_NVDLA_CSC_dl_for_check.scala 115:58:@46.4]
  wire  _T_257; // @[Mux.scala 46:19:@47.4]
  wire [5:0] _T_258; // @[Mux.scala 46:16:@48.4]
  wire  _T_259; // @[Mux.scala 46:19:@49.4]
  wire [6:0] pixel_x_init_w; // @[Mux.scala 46:16:@50.4]
  wire [6:0] pixel_x_init_offset_w; // @[NV_NVDLA_CSC_dl_for_check.scala 116:80:@52.4]
  wire [7:0] _T_264; // @[Cat.scala 30:58:@53.4]
  wire [6:0] _T_269; // @[Mux.scala 46:16:@56.4]
  wire [7:0] pixel_x_add_w; // @[Mux.scala 46:16:@58.4]
  wire [11:0] pixel_ch_stride_w; // @[Cat.scala 30:58:@59.4]
  wire [3:0] conv_y_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 126:74:@60.4]
  wire [5:0] _T_278; // @[NV_NVDLA_CSC_dl_for_check.scala 127:74:@63.4]
  wire [5:0] x_dilate_w; // @[NV_NVDLA_CSC_dl_for_check.scala 127:21:@64.4]
  wire [5:0] _T_282; // @[NV_NVDLA_CSC_dl_for_check.scala 128:74:@66.4]
  wire [5:0] y_dilate_w; // @[NV_NVDLA_CSC_dl_for_check.scala 128:21:@67.4]
  reg  layer_st_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 130:26:@68.4]
  reg [31:0] _RAND_0;
  reg [5:0] data_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 131:25:@70.4]
  reg [31:0] _RAND_1;
  reg [13:0] rls_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 132:25:@72.4]
  reg [31:0] _RAND_2;
  reg [13:0] h_offset_slice; // @[NV_NVDLA_CSC_dl_for_check.scala 133:29:@74.4]
  reg [31:0] _RAND_3;
  reg [16:0] entries; // @[NV_NVDLA_CSC_dl_for_check.scala 134:22:@76.4]
  reg [31:0] _RAND_4;
  reg [14:0] entries_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 135:28:@78.4]
  reg [31:0] _RAND_5;
  reg [12:0] dataout_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 136:32:@80.4]
  reg [31:0] _RAND_6;
  reg [28:0] rls_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 138:26:@84.4]
  reg [31:0] _RAND_7;
  reg [22:0] h_bias_0_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 139:30:@86.4]
  reg [31:0] _RAND_8;
  reg [30:0] h_bias_1_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 140:30:@88.4]
  reg [31:0] _RAND_9;
  reg [13:0] slice_left; // @[NV_NVDLA_CSC_dl_for_check.scala 141:25:@90.4]
  reg [31:0] _RAND_10;
  wire [14:0] entries_single_w; // @[NV_NVDLA_CSC_dl_for_check.scala 144:43:@91.4]
  wire [20:0] _T_353; // @[NV_NVDLA_CSC_dl_for_check.scala 145:41:@93.4]
  wire [14:0] entries_batch_w; // @[NV_NVDLA_CSC_dl_for_check.scala 145:56:@94.4]
  wire [16:0] entries_w; // @[NV_NVDLA_CSC_dl_for_check.scala 146:20:@97.4]
  wire [11:0] h_offset_slice_w; // @[NV_NVDLA_CSC_dl_for_check.scala 147:37:@98.4]
  wire [16:0] _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 148:33:@99.4]
  wire [22:0] h_bias_0_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 148:33:@99.4]
  wire [16:0] _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 149:33:@100.4]
  wire [30:0] h_bias_1_stride_w; // @[NV_NVDLA_CSC_dl_for_check.scala 149:33:@100.4]
  wire [12:0] rls_slices_w; // @[NV_NVDLA_CSC_dl_for_check.scala 150:41:@101.4]
  wire [13:0] _T_360; // @[NV_NVDLA_CSC_dl_for_check.scala 151:77:@102.4]
  wire [12:0] _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 151:113:@103.4]
  wire [13:0] _T_361; // @[NV_NVDLA_CSC_dl_for_check.scala 151:113:@103.4]
  wire [13:0] _T_362; // @[NV_NVDLA_CSC_dl_for_check.scala 151:113:@104.4]
  wire [13:0] slice_left_w; // @[NV_NVDLA_CSC_dl_for_check.scala 151:23:@105.4]
  wire [13:0] slices_oprand; // @[NV_NVDLA_CSC_dl_for_check.scala 152:24:@106.4]
  wire [14:0] _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 153:37:@107.4]
  wire [28:0] slice_entries_w; // @[NV_NVDLA_CSC_dl_for_check.scala 153:37:@107.4]
  reg [21:0] is_winograd_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 157:29:@111.4]
  reg [31:0] _RAND_11;
  reg [33:0] is_img_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 158:24:@113.4]
  reg [63:0] _RAND_12;
  reg [5:0] data_bank; // @[NV_NVDLA_CSC_dl_for_check.scala 159:24:@115.4]
  reg [31:0] _RAND_13;
  reg [13:0] datain_width; // @[NV_NVDLA_CSC_dl_for_check.scala 160:27:@117.4]
  reg [31:0] _RAND_14;
  reg [12:0] datain_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 161:31:@119.4]
  reg [31:0] _RAND_15;
  reg [12:0] datain_height_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 162:32:@121.4]
  reg [31:0] _RAND_16;
  reg [10:0] datain_channel_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 163:33:@123.4]
  reg [31:0] _RAND_17;
  reg [2:0] sub_h_total_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 164:29:@124.4]
  reg [31:0] _RAND_18;
  reg [2:0] sub_h_total_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 165:29:@125.4]
  reg [31:0] _RAND_19;
  reg [1:0] sub_h_total_g2; // @[NV_NVDLA_CSC_dl_for_check.scala 166:29:@126.4]
  reg [31:0] _RAND_20;
  reg [2:0] sub_h_total_g3; // @[NV_NVDLA_CSC_dl_for_check.scala 167:29:@127.4]
  reg [31:0] _RAND_21;
  reg [2:0] sub_h_total_g4; // @[NV_NVDLA_CSC_dl_for_check.scala 168:29:@128.4]
  reg [31:0] _RAND_22;
  reg [2:0] sub_h_total_g5; // @[NV_NVDLA_CSC_dl_for_check.scala 169:29:@129.4]
  reg [31:0] _RAND_23;
  reg [2:0] sub_h_total_g6; // @[NV_NVDLA_CSC_dl_for_check.scala 170:29:@130.4]
  reg [31:0] _RAND_24;
  reg [2:0] sub_h_total_g8; // @[NV_NVDLA_CSC_dl_for_check.scala 172:29:@132.4]
  reg [31:0] _RAND_25;
  reg [2:0] sub_h_total_g9; // @[NV_NVDLA_CSC_dl_for_check.scala 173:29:@133.4]
  reg [31:0] _RAND_26;
  reg [2:0] sub_h_total_g11; // @[NV_NVDLA_CSC_dl_for_check.scala 175:30:@135.4]
  reg [31:0] _RAND_27;
  reg [2:0] sub_h_cmp_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 176:27:@136.4]
  reg [31:0] _RAND_28;
  reg [2:0] sub_h_cmp_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 177:27:@137.4]
  reg [31:0] _RAND_29;
  reg [3:0] conv_x_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 178:28:@139.4]
  reg [31:0] _RAND_30;
  reg [3:0] conv_y_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 179:28:@141.4]
  reg [31:0] _RAND_31;
  reg [4:0] batch_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 181:24:@144.4]
  reg [31:0] _RAND_32;
  reg [6:0] pixel_x_init; // @[NV_NVDLA_CSC_dl_for_check.scala 182:27:@146.4]
  reg [31:0] _RAND_33;
  reg [6:0] pixel_x_init_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 183:34:@148.4]
  reg [31:0] _RAND_34;
  reg [7:0] pixel_x_add; // @[NV_NVDLA_CSC_dl_for_check.scala 184:26:@150.4]
  reg [31:0] _RAND_35;
  reg [6:0] pixel_x_byte_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 185:34:@152.4]
  reg [31:0] _RAND_36;
  reg [11:0] pixel_ch_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 186:30:@154.4]
  reg [31:0] _RAND_37;
  reg [5:0] x_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 187:23:@156.4]
  reg [31:0] _RAND_38;
  reg [5:0] y_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 188:23:@158.4]
  reg [31:0] _RAND_39;
  reg [15:0] pad_value; // @[NV_NVDLA_CSC_dl_for_check.scala 189:24:@160.4]
  reg [31:0] _RAND_40;
  reg [14:0] entries_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 190:26:@162.4]
  reg [31:0] _RAND_41;
  reg [16:0] h_bias_2_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 191:30:@164.4]
  reg [31:0] _RAND_42;
  reg [16:0] h_bias_3_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 192:30:@166.4]
  reg [31:0] _RAND_43;
  reg [13:0] last_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 194:26:@168.4]
  reg [31:0] _RAND_44;
  reg [28:0] last_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 195:27:@170.4]
  reg [31:0] _RAND_45;
  wire [33:0] _T_547; // @[Bitwise.scala 72:12:@178.6]
  wire [5:0] _T_549; // @[NV_NVDLA_CSC_dl_for_check.scala 202:38:@180.6]
  wire [13:0] _T_554; // @[NV_NVDLA_CSC_dl_for_check.scala 203:109:@184.6]
  wire [6:0] _T_557; // @[NV_NVDLA_CSC_dl_for_check.scala 206:109:@190.6]
  wire [10:0] _T_558; // @[NV_NVDLA_CSC_dl_for_check.scala 206:30:@191.6]
  wire [1:0] _T_559; // @[NV_NVDLA_CSC_dl_for_check.scala 209:36:@195.6]
  wire [14:0] _T_562; // @[Cat.scala 30:58:@224.6]
  wire [21:0] _GEN_0; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [33:0] _GEN_1; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [5:0] _GEN_2; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [13:0] _GEN_3; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [12:0] _GEN_4; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [12:0] _GEN_5; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [10:0] _GEN_6; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_7; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_8; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [1:0] _GEN_9; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_10; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_11; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_12; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_13; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_15; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_16; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_18; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_19; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [2:0] _GEN_20; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [3:0] _GEN_21; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [3:0] _GEN_22; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [5:0] _GEN_24; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [4:0] _GEN_25; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [6:0] _GEN_26; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [6:0] _GEN_27; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [7:0] _GEN_28; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [6:0] _GEN_29; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [11:0] _GEN_30; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [5:0] _GEN_31; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [5:0] _GEN_32; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [15:0] _GEN_33; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [16:0] _GEN_34; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [14:0] _GEN_35; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [14:0] _GEN_36; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [13:0] _GEN_37; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [13:0] _GEN_38; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [13:0] _GEN_39; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [12:0] _GEN_40; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  wire [22:0] _GEN_43; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  wire [30:0] _GEN_44; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  wire [16:0] _GEN_45; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  wire [16:0] _GEN_46; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  wire [28:0] _GEN_47; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  wire [13:0] _GEN_48; // @[NV_NVDLA_CSC_dl_for_check.scala 251:17:@244.4]
  wire [28:0] _GEN_49; // @[NV_NVDLA_CSC_dl_for_check.scala 251:17:@244.4]
  reg [14:0] dat_entry_st; // @[NV_NVDLA_CSC_dl_for_check.scala 274:59:@269.4]
  reg [31:0] _RAND_46;
  wire  _T_643; // @[NV_NVDLA_CSC_dl_for_check.scala 315:37:@328.4]
  wire  _T_644; // @[NV_NVDLA_CSC_dl_for_check.scala 315:23:@329.4]
  wire  _T_1517; // @[NV_NVDLA_CSC_dl_for_check.scala 911:32:@1247.4]
  reg  dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 896:41:@1215.4]
  reg [31:0] _RAND_47;
  wire  _T_1518; // @[NV_NVDLA_CSC_dl_for_check.scala 911:36:@1248.4]
  wire  _T_1519; // @[NV_NVDLA_CSC_dl_for_check.scala 912:35:@1249.4]
  reg  dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 896:41:@1213.4]
  reg [31:0] _RAND_48;
  wire  _T_1520; // @[NV_NVDLA_CSC_dl_for_check.scala 912:39:@1250.4]
  wire  _T_1521; // @[NV_NVDLA_CSC_dl_for_check.scala 911:57:@1251.4]
  wire  _T_1522; // @[NV_NVDLA_CSC_dl_for_check.scala 913:35:@1252.4]
  reg  dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 896:41:@1212.4]
  reg [31:0] _RAND_49;
  wire  _T_1523; // @[NV_NVDLA_CSC_dl_for_check.scala 913:39:@1253.4]
  wire  dat_rsp_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 912:60:@1254.4]
  wire  _T_1525; // @[NV_NVDLA_CSC_dl_for_check.scala 920:42:@1256.4]
  wire [26:0] _T_1529; // @[Bitwise.scala 72:12:@1258.4]
  reg [26:0] _T_1507; // @[NV_NVDLA_CSC_dl_for_check.scala 898:41:@1220.4]
  reg [31:0] _RAND_50;
  wire [26:0] _T_1530; // @[NV_NVDLA_CSC_dl_for_check.scala 920:47:@1259.4]
  wire  _T_1531; // @[NV_NVDLA_CSC_dl_for_check.scala 921:42:@1260.4]
  wire [26:0] _T_1535; // @[Bitwise.scala 72:12:@1262.4]
  reg [26:0] _T_1501; // @[NV_NVDLA_CSC_dl_for_check.scala 898:41:@1218.4]
  reg [31:0] _RAND_51;
  wire [26:0] _T_1536; // @[NV_NVDLA_CSC_dl_for_check.scala 921:47:@1263.4]
  wire [26:0] _T_1537; // @[NV_NVDLA_CSC_dl_for_check.scala 920:66:@1264.4]
  wire  _T_1538; // @[NV_NVDLA_CSC_dl_for_check.scala 922:42:@1265.4]
  wire [26:0] _T_1542; // @[Bitwise.scala 72:12:@1267.4]
  reg [26:0] _T_1498; // @[NV_NVDLA_CSC_dl_for_check.scala 898:41:@1217.4]
  reg [31:0] _RAND_52;
  wire [26:0] _T_1543; // @[NV_NVDLA_CSC_dl_for_check.scala 922:47:@1268.4]
  wire [26:0] dat_rsp_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 921:66:@1269.4]
  wire  dat_rsp_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 946:26:@1288.4]
  wire  sub_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 312:29:@327.4]
  wire  _T_646; // @[NV_NVDLA_CSC_dl_for_check.scala 315:66:@330.4]
  wire  _T_647; // @[NV_NVDLA_CSC_dl_for_check.scala 315:53:@331.4]
  wire  dat_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 315:42:@332.4]
  wire [13:0] sc2cdma_dat_slices_w; // @[NV_NVDLA_CSC_dl_for_check.scala 316:28:@334.4]
  wire [28:0] _T_650; // @[NV_NVDLA_CSC_dl_for_check.scala 317:29:@336.4]
  wire [14:0] sc2cdma_dat_entries_w; // @[NV_NVDLA_CSC_dl_for_check.scala 271:34:@266.4 NV_NVDLA_CSC_dl_for_check.scala 317:23:@337.4]
  wire [14:0] dat_entry_avl_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 284:28:@278.4]
  wire [15:0] _T_600; // @[NV_NVDLA_CSC_dl_for_check.scala 289:37:@283.4]
  wire [14:0] dat_entry_st_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 289:37:@284.4]
  wire [14:0] _T_606; // @[Cat.scala 30:58:@286.4]
  wire [15:0] _T_607; // @[NV_NVDLA_CSC_dl_for_check.scala 290:46:@287.4]
  wire [15:0] _T_608; // @[NV_NVDLA_CSC_dl_for_check.scala 290:46:@288.4]
  wire [14:0] dat_entry_st_inc_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 290:46:@289.4]
  wire  is_dat_entry_st_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 291:45:@292.4]
  wire [14:0] _T_616; // @[NV_NVDLA_CSC_dl_for_check.scala 292:83:@293.4]
  wire [14:0] dat_entry_st_w; // @[NV_NVDLA_CSC_dl_for_check.scala 292:25:@294.4]
  wire  _T_638; // @[NV_NVDLA_CSC_dl_for_check.scala 303:13:@317.4]
  wire [14:0] _GEN_55; // @[NV_NVDLA_CSC_dl_for_check.scala 303:25:@318.4]
  reg  _T_653; // @[NV_NVDLA_CSC_dl_for_check.scala 319:37:@338.4]
  reg [31:0] _RAND_53;
  reg [13:0] _T_656; // @[Reg.scala 19:20:@341.4]
  reg [31:0] _RAND_54;
  wire [13:0] _GEN_57; // @[Reg.scala 20:19:@342.4]
  reg [14:0] _T_659; // @[Reg.scala 19:20:@346.4]
  reg [31:0] _RAND_55;
  wire [14:0] _GEN_58; // @[Reg.scala 20:19:@347.4]
  reg  _T_664; // @[NV_NVDLA_CSC_dl_for_check.scala 333:50:@352.4]
  reg [31:0] _RAND_56;
  reg  _T_667; // @[NV_NVDLA_CSC_dl_for_check.scala 333:50:@353.4]
  reg [31:0] _RAND_57;
  reg  _T_670; // @[NV_NVDLA_CSC_dl_for_check.scala 333:50:@354.4]
  reg [31:0] _RAND_58;
  reg  _T_673; // @[NV_NVDLA_CSC_dl_for_check.scala 333:50:@355.4]
  reg [31:0] _RAND_59;
  reg  _T_676; // @[NV_NVDLA_CSC_dl_for_check.scala 333:50:@356.4]
  reg [31:0] _RAND_60;
  reg [30:0] _T_681; // @[NV_NVDLA_CSC_dl_for_check.scala 335:47:@358.4]
  reg [31:0] _RAND_61;
  reg [30:0] _T_684; // @[NV_NVDLA_CSC_dl_for_check.scala 335:47:@359.4]
  reg [31:0] _RAND_62;
  reg [30:0] _T_687; // @[NV_NVDLA_CSC_dl_for_check.scala 335:47:@360.4]
  reg [31:0] _RAND_63;
  reg [30:0] _T_690; // @[NV_NVDLA_CSC_dl_for_check.scala 335:47:@361.4]
  reg [31:0] _RAND_64;
  reg [30:0] _T_693; // @[NV_NVDLA_CSC_dl_for_check.scala 335:47:@362.4]
  reg [31:0] _RAND_65;
  wire [30:0] _GEN_59; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@366.4]
  wire [30:0] _GEN_60; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@370.4]
  wire [30:0] _GEN_61; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@374.4]
  wire [30:0] _GEN_62; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@378.4]
  wire [30:0] _GEN_63; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@382.4]
  wire  _T_694; // @[NV_NVDLA_CSC_dl_for_check.scala 347:36:@385.4]
  wire  dl_in_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 347:21:@386.4]
  wire  _T_695; // @[NV_NVDLA_CSC_dl_for_check.scala 348:34:@387.4]
  wire [30:0] dl_in_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 348:19:@388.4]
  reg  _T_700; // @[NV_NVDLA_CSC_dl_for_check.scala 352:36:@390.4]
  reg [31:0] _RAND_66;
  reg  _T_703; // @[NV_NVDLA_CSC_dl_for_check.scala 352:36:@391.4]
  reg [31:0] _RAND_67;
  reg  _T_706; // @[NV_NVDLA_CSC_dl_for_check.scala 352:36:@392.4]
  reg [31:0] _RAND_68;
  reg  _T_709; // @[NV_NVDLA_CSC_dl_for_check.scala 352:36:@393.4]
  reg [31:0] _RAND_69;
  reg [30:0] _T_714; // @[NV_NVDLA_CSC_dl_for_check.scala 354:34:@395.4]
  reg [31:0] _RAND_70;
  reg [30:0] _T_717; // @[NV_NVDLA_CSC_dl_for_check.scala 354:34:@396.4]
  reg [31:0] _RAND_71;
  reg [30:0] _T_720; // @[NV_NVDLA_CSC_dl_for_check.scala 354:34:@397.4]
  reg [31:0] _RAND_72;
  reg [30:0] _T_723; // @[NV_NVDLA_CSC_dl_for_check.scala 354:34:@398.4]
  reg [31:0] _RAND_73;
  wire [30:0] _GEN_64; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@402.4]
  wire [30:0] _GEN_65; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@406.4]
  wire [30:0] _GEN_66; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@410.4]
  wire [30:0] _GEN_67; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@414.4]
  wire  _T_724; // @[NV_NVDLA_CSC_dl_for_check.scala 366:30:@417.4]
  wire  _T_725; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@418.4]
  wire  _T_726; // @[NV_NVDLA_CSC_dl_for_check.scala 367:30:@419.4]
  wire  _T_727; // @[NV_NVDLA_CSC_dl_for_check.scala 367:34:@420.4]
  wire  _T_728; // @[NV_NVDLA_CSC_dl_for_check.scala 366:50:@421.4]
  wire  _T_729; // @[NV_NVDLA_CSC_dl_for_check.scala 368:30:@422.4]
  wire  _T_730; // @[NV_NVDLA_CSC_dl_for_check.scala 368:34:@423.4]
  wire  dl_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 367:50:@424.4]
  wire  _T_731; // @[NV_NVDLA_CSC_dl_for_check.scala 370:37:@425.4]
  wire [30:0] _T_735; // @[Bitwise.scala 72:12:@427.4]
  wire [30:0] _T_736; // @[NV_NVDLA_CSC_dl_for_check.scala 370:42:@428.4]
  wire  _T_737; // @[NV_NVDLA_CSC_dl_for_check.scala 371:37:@429.4]
  wire [30:0] _T_741; // @[Bitwise.scala 72:12:@431.4]
  wire [30:0] _T_742; // @[NV_NVDLA_CSC_dl_for_check.scala 371:42:@432.4]
  wire [30:0] _T_743; // @[NV_NVDLA_CSC_dl_for_check.scala 370:56:@433.4]
  wire  _T_744; // @[NV_NVDLA_CSC_dl_for_check.scala 372:37:@434.4]
  wire [30:0] _T_748; // @[Bitwise.scala 72:12:@436.4]
  wire [30:0] _T_749; // @[NV_NVDLA_CSC_dl_for_check.scala 372:42:@437.4]
  wire [30:0] dl_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 371:56:@438.4]
  wire [4:0] dl_w_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 375:24:@439.4]
  wire [4:0] dl_h_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 376:24:@440.4]
  wire [6:0] dl_channel_size; // @[NV_NVDLA_CSC_dl_for_check.scala 377:28:@441.4]
  wire [6:0] dl_stripe_length; // @[NV_NVDLA_CSC_dl_for_check.scala 378:29:@442.4]
  wire [1:0] dl_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 379:25:@443.4]
  wire  dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 380:25:@444.4]
  wire  dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 381:27:@445.4]
  wire  dl_group_end; // @[NV_NVDLA_CSC_dl_for_check.scala 382:25:@446.4]
  wire  dl_layer_end; // @[NV_NVDLA_CSC_dl_for_check.scala 383:25:@447.4]
  wire  dl_dat_release; // @[NV_NVDLA_CSC_dl_for_check.scala 384:27:@448.4]
  reg [4:0] batch_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 389:24:@451.4]
  reg [31:0] _RAND_74;
  reg [6:0] stripe_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 412:25:@476.4]
  reg [31:0] _RAND_75;
  wire  _T_806; // @[NV_NVDLA_CSC_dl_for_check.scala 439:37:@505.4]
  wire  _T_807; // @[NV_NVDLA_CSC_dl_for_check.scala 439:24:@506.4]
  reg [1:0] sub_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 401:24:@461.4]
  reg [31:0] _RAND_76;
  wire  _T_809; // @[NV_NVDLA_CSC_dl_for_check.scala 439:56:@507.4]
  wire  _T_810; // @[NV_NVDLA_CSC_dl_for_check.scala 439:44:@508.4]
  wire  _T_811; // @[NV_NVDLA_CSC_dl_for_check.scala 439:42:@509.4]
  wire  _T_813; // @[NV_NVDLA_CSC_dl_for_check.scala 439:75:@510.4]
  wire  _T_814; // @[NV_NVDLA_CSC_dl_for_check.scala 439:63:@511.4]
  wire  _T_815; // @[NV_NVDLA_CSC_dl_for_check.scala 439:61:@512.4]
  reg  dat_exec_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 431:32:@498.4]
  reg [31:0] _RAND_77;
  wire  _T_817; // @[NV_NVDLA_CSC_dl_for_check.scala 439:22:@513.4]
  wire  dat_exec_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 438:22:@514.4]
  wire  _T_754; // @[NV_NVDLA_CSC_dl_for_check.scala 391:15:@452.4]
  wire [5:0] _T_758; // @[NV_NVDLA_CSC_dl_for_check.scala 394:28:@454.6]
  wire  is_batch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 398:27:@459.4]
  wire [5:0] _T_759; // @[NV_NVDLA_CSC_dl_for_check.scala 393:21:@455.6]
  wire [5:0] _T_760; // @[NV_NVDLA_CSC_dl_for_check.scala 392:21:@456.6]
  wire [5:0] _GEN_68; // @[NV_NVDLA_CSC_dl_for_check.scala 391:32:@453.4]
  wire [2:0] sub_h_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 404:31:@463.4]
  wire  is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 405:32:@464.4]
  wire  _T_767; // @[NV_NVDLA_CSC_dl_for_check.scala 406:51:@466.4]
  wire  _T_769; // @[NV_NVDLA_CSC_dl_for_check.scala 406:82:@467.4]
  wire  _T_770; // @[NV_NVDLA_CSC_dl_for_check.scala 406:55:@468.4]
  wire  _T_771; // @[NV_NVDLA_CSC_dl_for_check.scala 406:88:@469.4]
  wire  sub_h_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 406:33:@470.4]
  wire  _T_772; // @[NV_NVDLA_CSC_dl_for_check.scala 408:31:@472.6]
  wire [2:0] _T_774; // @[NV_NVDLA_CSC_dl_for_check.scala 408:21:@473.6]
  wire [2:0] _GEN_69; // @[NV_NVDLA_CSC_dl_for_check.scala 407:23:@471.4]
  wire [7:0] _T_780; // @[NV_NVDLA_CSC_dl_for_check.scala 416:34:@479.4]
  wire [6:0] stripe_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 416:41:@480.4]
  wire  _T_781; // @[NV_NVDLA_CSC_dl_for_check.scala 417:51:@481.4]
  wire  is_stripe_equal; // @[NV_NVDLA_CSC_dl_for_check.scala 417:33:@482.4]
  wire  is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 418:34:@484.4]
  wire  _T_784; // @[NV_NVDLA_CSC_dl_for_check.scala 419:52:@486.4]
  wire  stripe_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 419:34:@487.4]
  wire  _T_786; // @[NV_NVDLA_CSC_dl_for_check.scala 423:41:@489.6]
  wire  _T_787; // @[NV_NVDLA_CSC_dl_for_check.scala 423:39:@490.6]
  wire [6:0] _T_789; // @[NV_NVDLA_CSC_dl_for_check.scala 424:22:@491.6]
  wire [6:0] _T_790; // @[NV_NVDLA_CSC_dl_for_check.scala 423:22:@492.6]
  wire [6:0] _T_791; // @[NV_NVDLA_CSC_dl_for_check.scala 422:22:@493.6]
  wire [6:0] _GEN_70; // @[NV_NVDLA_CSC_dl_for_check.scala 421:24:@488.4]
  reg  dat_pipe_local_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 429:35:@496.4]
  reg [31:0] _RAND_78;
  reg  dat_pipe_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 430:32:@497.4]
  reg [31:0] _RAND_79;
  wire  dat_pipe_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 437:27:@503.4]
  wire  _T_799; // @[NV_NVDLA_CSC_dl_for_check.scala 434:49:@500.4]
  wire  _T_802; // @[NV_NVDLA_CSC_dl_for_check.scala 435:32:@501.4]
  wire  dat_pipe_local_valid_w; // @[NV_NVDLA_CSC_dl_for_check.scala 434:33:@502.4]
  reg [7:0] dat_req_bytes_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 447:31:@519.4]
  reg [31:0] _RAND_80;
  wire [7:0] dat_req_bytes; // @[Cat.scala 30:58:@520.4]
  wire [7:0] _GEN_71; // @[NV_NVDLA_CSC_dl_for_check.scala 449:21:@521.4]
  reg [12:0] dataout_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 455:28:@524.4]
  reg [31:0] _RAND_81;
  reg [12:0] dataout_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 456:28:@525.4]
  reg [31:0] _RAND_82;
  wire [12:0] _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 459:39:@526.4]
  wire [13:0] _T_826; // @[NV_NVDLA_CSC_dl_for_check.scala 459:39:@526.4]
  wire [12:0] dataout_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 459:39:@527.4]
  wire  _T_827; // @[NV_NVDLA_CSC_dl_for_check.scala 460:29:@528.4]
  wire  _T_828; // @[NV_NVDLA_CSC_dl_for_check.scala 460:61:@529.4]
  wire  is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 460:44:@530.4]
  wire  _T_830; // @[NV_NVDLA_CSC_dl_for_check.scala 463:43:@533.4]
  wire  _T_831; // @[NV_NVDLA_CSC_dl_for_check.scala 463:41:@534.4]
  wire [12:0] _T_832; // @[NV_NVDLA_CSC_dl_for_check.scala 464:26:@535.4]
  wire [12:0] _T_833; // @[NV_NVDLA_CSC_dl_for_check.scala 463:26:@536.4]
  wire [12:0] dataout_w_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 462:26:@537.4]
  wire  _T_835; // @[NV_NVDLA_CSC_dl_for_check.scala 465:70:@539.4]
  wire  dataout_w_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 465:37:@540.4]
  wire  _T_836; // @[NV_NVDLA_CSC_dl_for_check.scala 466:55:@541.4]
  wire  _T_837; // @[NV_NVDLA_CSC_dl_for_check.scala 466:71:@542.4]
  wire  dataout_w_ori_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 466:37:@543.4]
  wire [12:0] _GEN_72; // @[NV_NVDLA_CSC_dl_for_check.scala 468:27:@544.4]
  wire [12:0] _GEN_73; // @[NV_NVDLA_CSC_dl_for_check.scala 471:27:@547.4]
  reg [10:0] datain_c_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 476:27:@550.4]
  reg [31:0] _RAND_83;
  wire  is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 478:37:@551.4]
  wire  _T_841; // @[NV_NVDLA_CSC_dl_for_check.scala 479:70:@553.4]
  wire  datain_c_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 479:36:@554.4]
  wire [11:0] _T_845; // @[NV_NVDLA_CSC_dl_for_check.scala 484:34:@556.6]
  wire [10:0] _T_846; // @[NV_NVDLA_CSC_dl_for_check.scala 484:34:@557.6]
  wire [10:0] _T_847; // @[NV_NVDLA_CSC_dl_for_check.scala 483:24:@558.6]
  wire [10:0] _T_848; // @[NV_NVDLA_CSC_dl_for_check.scala 482:24:@559.6]
  wire [10:0] _GEN_74; // @[NV_NVDLA_CSC_dl_for_check.scala 481:26:@555.4]
  reg [13:0] datain_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 488:27:@562.4]
  reg [31:0] _RAND_84;
  reg [13:0] datain_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 489:27:@563.4]
  reg [31:0] _RAND_85;
  reg [15:0] pixel_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 490:26:@564.4]
  reg [31:0] _RAND_86;
  reg [15:0] pixel_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 491:26:@565.4]
  reg [31:0] _RAND_87;
  reg [15:0] pixel_w_ch_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 492:29:@566.4]
  reg [31:0] _RAND_88;
  reg [12:0] channel_op_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 493:29:@567.4]
  reg [31:0] _RAND_89;
  reg  pixel_force_clr_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 495:33:@569.4]
  reg [31:0] _RAND_90;
  reg  pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 496:35:@570.4]
  reg [31:0] _RAND_91;
  wire [12:0] _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 500:41:@571.4]
  wire [13:0] _T_869; // @[NV_NVDLA_CSC_dl_for_check.scala 500:41:@571.4]
  wire [13:0] _T_870; // @[NV_NVDLA_CSC_dl_for_check.scala 500:41:@572.4]
  wire [13:0] datain_w_cnt_st; // @[NV_NVDLA_CSC_dl_for_check.scala 498:26:@574.4]
  wire  _T_872; // @[NV_NVDLA_CSC_dl_for_check.scala 501:42:@575.4]
  wire [14:0] _T_874; // @[NV_NVDLA_CSC_dl_for_check.scala 501:60:@576.4]
  wire [13:0] _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 501:81:@577.4]
  wire [14:0] _T_875; // @[NV_NVDLA_CSC_dl_for_check.scala 501:81:@577.4]
  wire [14:0] datain_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 501:27:@578.4]
  wire [14:0] _T_878; // @[NV_NVDLA_CSC_dl_for_check.scala 506:25:@581.4]
  wire [14:0] _T_879; // @[NV_NVDLA_CSC_dl_for_check.scala 505:25:@582.4]
  wire [14:0] datain_w_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 504:25:@583.4]
  wire [5:0] _GEN_693; // @[NV_NVDLA_CSC_dl_for_check.scala 508:35:@584.4]
  wire [10:0] dl_w_offset_ext; // @[NV_NVDLA_CSC_dl_for_check.scala 508:35:@584.4]
  wire [13:0] _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 509:34:@585.4]
  wire [14:0] _T_880; // @[NV_NVDLA_CSC_dl_for_check.scala 509:34:@585.4]
  wire [13:0] datain_w_cur; // @[NV_NVDLA_CSC_dl_for_check.scala 509:53:@586.4]
  wire  _T_883; // @[NV_NVDLA_CSC_dl_for_check.scala 510:96:@589.4]
  wire  _T_884; // @[NV_NVDLA_CSC_dl_for_check.scala 510:86:@590.4]
  wire  _T_885; // @[NV_NVDLA_CSC_dl_for_check.scala 510:84:@591.4]
  wire  datain_w_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 510:36:@592.4]
  wire  _T_888; // @[NV_NVDLA_CSC_dl_for_check.scala 511:99:@595.4]
  wire  _T_889; // @[NV_NVDLA_CSC_dl_for_check.scala 511:89:@596.4]
  wire  _T_890; // @[NV_NVDLA_CSC_dl_for_check.scala 511:87:@597.4]
  wire  datain_w_ori_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 511:36:@598.4]
  wire [7:0] pixel_x_cnt_add; // @[NV_NVDLA_CSC_dl_for_check.scala 514:26:@599.4]
  wire  _T_894; // @[NV_NVDLA_CSC_dl_for_check.scala 516:79:@601.4]
  wire [7:0] _T_898; // @[NV_NVDLA_CSC_dl_for_check.scala 517:75:@604.4]
  wire [7:0] total_channel_op; // @[NV_NVDLA_CSC_dl_for_check.scala 516:27:@605.4]
  wire  _T_899; // @[NV_NVDLA_CSC_dl_for_check.scala 518:37:@606.4]
  wire  _T_901; // @[NV_NVDLA_CSC_dl_for_check.scala 519:35:@607.4]
  wire [13:0] _T_903; // @[NV_NVDLA_CSC_dl_for_check.scala 519:66:@608.4]
  wire [13:0] _T_904; // @[NV_NVDLA_CSC_dl_for_check.scala 519:22:@609.4]
  wire [13:0] _T_905; // @[NV_NVDLA_CSC_dl_for_check.scala 518:22:@610.4]
  wire [12:0] _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 521:44:@612.4]
  wire  next_is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 521:44:@612.4]
  wire  _T_906; // @[NV_NVDLA_CSC_dl_for_check.scala 525:39:@613.4]
  wire  _T_907; // @[NV_NVDLA_CSC_dl_for_check.scala 525:54:@614.4]
  wire  _T_908; // @[NV_NVDLA_CSC_dl_for_check.scala 525:71:@615.4]
  wire  _T_911; // @[NV_NVDLA_CSC_dl_for_check.scala 526:73:@618.4]
  wire  _T_912; // @[NV_NVDLA_CSC_dl_for_check.scala 526:71:@619.4]
  wire [15:0] _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 526:99:@620.4]
  wire [16:0] _T_913; // @[NV_NVDLA_CSC_dl_for_check.scala 526:99:@620.4]
  wire  _T_915; // @[NV_NVDLA_CSC_dl_for_check.scala 527:54:@622.4]
  wire [15:0] _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 527:90:@623.4]
  wire [16:0] _T_916; // @[NV_NVDLA_CSC_dl_for_check.scala 527:90:@623.4]
  wire  _T_918; // @[NV_NVDLA_CSC_dl_for_check.scala 528:56:@625.4]
  wire  _T_919; // @[NV_NVDLA_CSC_dl_for_check.scala 528:54:@626.4]
  wire [16:0] _T_921; // @[NV_NVDLA_CSC_dl_for_check.scala 528:91:@627.4]
  wire  _T_922; // @[NV_NVDLA_CSC_dl_for_check.scala 529:41:@628.4]
  wire  _T_923; // @[NV_NVDLA_CSC_dl_for_check.scala 529:39:@629.4]
  wire [15:0] _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 529:81:@630.4]
  wire [16:0] _T_924; // @[NV_NVDLA_CSC_dl_for_check.scala 529:81:@630.4]
  wire [16:0] _T_925; // @[NV_NVDLA_CSC_dl_for_check.scala 529:24:@631.4]
  wire [16:0] _T_926; // @[NV_NVDLA_CSC_dl_for_check.scala 528:24:@632.4]
  wire [16:0] _T_927; // @[NV_NVDLA_CSC_dl_for_check.scala 527:24:@633.4]
  wire [16:0] _T_928; // @[NV_NVDLA_CSC_dl_for_check.scala 526:24:@634.4]
  wire [16:0] _T_929; // @[NV_NVDLA_CSC_dl_for_check.scala 525:24:@635.4]
  wire [16:0] pixel_w_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 524:24:@636.4]
  wire [9:0] _T_935; // @[NV_NVDLA_CSC_dl_for_check.scala 531:68:@638.4]
  wire [14:0] pixel_w_cur; // @[Cat.scala 30:58:@639.4]
  wire  _T_944; // @[NV_NVDLA_CSC_dl_for_check.scala 534:68:@650.4]
  wire  _T_945; // @[NV_NVDLA_CSC_dl_for_check.scala 534:57:@651.4]
  wire  _T_946; // @[NV_NVDLA_CSC_dl_for_check.scala 534:72:@652.4]
  wire  _T_947; // @[NV_NVDLA_CSC_dl_for_check.scala 534:88:@653.4]
  wire  _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 534:103:@654.4]
  wire  pixel_ch_ori_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 534:39:@655.4]
  wire  _T_950; // @[NV_NVDLA_CSC_dl_for_check.scala 536:42:@657.4]
  wire  _T_953; // @[NV_NVDLA_CSC_dl_for_check.scala 536:74:@658.4]
  wire  pixel_force_fetch; // @[NV_NVDLA_CSC_dl_for_check.scala 536:28:@659.4]
  wire  _T_955; // @[NV_NVDLA_CSC_dl_for_check.scala 537:36:@661.4]
  wire  _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 537:72:@662.4]
  wire  pixel_force_clr; // @[NV_NVDLA_CSC_dl_for_check.scala 537:51:@663.4]
  wire [14:0] _GEN_75; // @[NV_NVDLA_CSC_dl_for_check.scala 539:26:@664.4]
  wire [16:0] _GEN_76; // @[NV_NVDLA_CSC_dl_for_check.scala 539:26:@664.4]
  wire [14:0] _GEN_77; // @[NV_NVDLA_CSC_dl_for_check.scala 543:26:@668.4]
  wire [16:0] _GEN_78; // @[NV_NVDLA_CSC_dl_for_check.scala 543:26:@668.4]
  wire [16:0] _GEN_79; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@672.4]
  reg [13:0] datain_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 553:27:@675.4]
  reg [31:0] _RAND_92;
  reg [13:0] datain_h_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 554:27:@676.4]
  reg [31:0] _RAND_93;
  wire [13:0] _GEN_699; // @[NV_NVDLA_CSC_dl_for_check.scala 556:77:@677.4]
  wire [14:0] _T_963; // @[NV_NVDLA_CSC_dl_for_check.scala 556:77:@677.4]
  wire [14:0] datain_h_cnt_st; // @[NV_NVDLA_CSC_dl_for_check.scala 556:77:@678.4]
  wire [13:0] _GEN_700; // @[NV_NVDLA_CSC_dl_for_check.scala 557:37:@680.4]
  wire [14:0] _T_965; // @[NV_NVDLA_CSC_dl_for_check.scala 557:37:@680.4]
  wire [13:0] datain_h_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 557:37:@681.4]
  wire  _T_966; // @[NV_NVDLA_CSC_dl_for_check.scala 558:52:@682.4]
  wire  _T_967; // @[NV_NVDLA_CSC_dl_for_check.scala 558:35:@683.4]
  wire [13:0] _T_970; // @[NV_NVDLA_CSC_dl_for_check.scala 560:25:@686.4]
  wire [13:0] _T_971; // @[NV_NVDLA_CSC_dl_for_check.scala 559:25:@687.4]
  wire [14:0] datain_h_cnt_w; // @[NV_NVDLA_CSC_dl_for_check.scala 558:25:@688.4]
  wire  _T_974; // @[NV_NVDLA_CSC_dl_for_check.scala 561:91:@691.4]
  wire  _T_975; // @[NV_NVDLA_CSC_dl_for_check.scala 561:54:@692.4]
  wire  datain_h_cnt_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 561:36:@693.4]
  wire [5:0] _GEN_701; // @[NV_NVDLA_CSC_dl_for_check.scala 563:35:@697.4]
  wire [10:0] dl_h_offset_ext; // @[NV_NVDLA_CSC_dl_for_check.scala 563:35:@697.4]
  wire [13:0] _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 564:34:@698.4]
  wire [14:0] _T_978; // @[NV_NVDLA_CSC_dl_for_check.scala 564:34:@698.4]
  wire [14:0] _GEN_703; // @[NV_NVDLA_CSC_dl_for_check.scala 564:53:@699.4]
  wire [15:0] _T_979; // @[NV_NVDLA_CSC_dl_for_check.scala 564:53:@699.4]
  wire [13:0] datain_h_cur; // @[NV_NVDLA_CSC_dl_for_check.scala 564:66:@700.4]
  wire [14:0] _GEN_80; // @[NV_NVDLA_CSC_dl_for_check.scala 566:26:@701.4]
  wire [14:0] _GEN_81; // @[NV_NVDLA_CSC_dl_for_check.scala 567:26:@704.4]
  wire  _T_980; // @[NV_NVDLA_CSC_dl_for_check.scala 570:39:@707.4]
  wire [13:0] _GEN_704; // @[NV_NVDLA_CSC_dl_for_check.scala 570:59:@708.4]
  wire  _T_981; // @[NV_NVDLA_CSC_dl_for_check.scala 570:59:@708.4]
  wire  _T_982; // @[NV_NVDLA_CSC_dl_for_check.scala 570:44:@709.4]
  wire  _T_983; // @[NV_NVDLA_CSC_dl_for_check.scala 570:92:@710.4]
  wire  _T_984; // @[NV_NVDLA_CSC_dl_for_check.scala 570:78:@711.4]
  wire [13:0] _GEN_705; // @[NV_NVDLA_CSC_dl_for_check.scala 570:112:@712.4]
  wire  _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 570:112:@712.4]
  wire  dat_conv_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 570:97:@713.4]
  wire [11:0] _T_986; // @[NV_NVDLA_CSC_dl_for_check.scala 572:35:@714.4]
  wire  _T_988; // @[NV_NVDLA_CSC_dl_for_check.scala 572:43:@715.4]
  wire  _T_989; // @[NV_NVDLA_CSC_dl_for_check.scala 572:61:@716.4]
  wire  _T_990; // @[NV_NVDLA_CSC_dl_for_check.scala 572:47:@717.4]
  wire [5:0] _T_991; // @[NV_NVDLA_CSC_dl_for_check.scala 572:77:@718.4]
  wire  _T_993; // @[NV_NVDLA_CSC_dl_for_check.scala 572:84:@719.4]
  wire  dat_wg_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 572:65:@720.4]
  wire  dat_img_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 573:42:@723.4]
  wire  _T_1080; // @[NV_NVDLA_CSC_dl_for_check.scala 659:33:@821.4]
  wire  _T_1081; // @[NV_NVDLA_CSC_dl_for_check.scala 660:38:@822.4]
  wire  _T_1082; // @[NV_NVDLA_CSC_dl_for_check.scala 661:24:@823.4]
  wire  _T_1084; // @[NV_NVDLA_CSC_dl_for_check.scala 661:41:@825.4]
  wire [12:0] _T_1086; // @[NV_NVDLA_CSC_dl_for_check.scala 661:97:@826.4]
  wire [14:0] _T_1087; // @[Cat.scala 30:58:@827.4]
  wire  _T_1089; // @[NV_NVDLA_CSC_dl_for_check.scala 662:38:@828.4]
  wire [11:0] _T_1094; // @[NV_NVDLA_CSC_dl_for_check.scala 663:54:@831.4]
  wire [14:0] _T_1095; // @[Cat.scala 30:58:@832.4]
  wire [14:0] _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 662:23:@833.4]
  wire [14:0] _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 661:23:@834.4]
  wire [14:0] _T_1098; // @[NV_NVDLA_CSC_dl_for_check.scala 660:23:@835.4]
  wire [14:0] w_bias_int8; // @[NV_NVDLA_CSC_dl_for_check.scala 659:23:@836.4]
  wire [13:0] w_bias_w; // @[NV_NVDLA_CSC_dl_for_check.scala 673:24:@838.4]
  wire [11:0] _T_997; // @[NV_NVDLA_CSC_dl_for_check.scala 577:32:@725.4]
  wire [14:0] _GEN_707; // @[NV_NVDLA_CSC_dl_for_check.scala 577:40:@726.4]
  wire  dat_img_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 577:40:@726.4]
  wire  _T_998; // @[NV_NVDLA_CSC_dl_for_check.scala 578:34:@727.4]
  wire  _T_999; // @[NV_NVDLA_CSC_dl_for_check.scala 578:76:@728.4]
  wire  _T_1000; // @[NV_NVDLA_CSC_dl_for_check.scala 578:61:@729.4]
  wire  dat_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 578:24:@730.4]
  wire  _T_1001; // @[NV_NVDLA_CSC_dl_for_check.scala 579:35:@731.4]
  wire  _T_1002; // @[NV_NVDLA_CSC_dl_for_check.scala 579:39:@732.4]
  wire  _T_1003; // @[NV_NVDLA_CSC_dl_for_check.scala 579:70:@733.4]
  wire  _T_1004; // @[NV_NVDLA_CSC_dl_for_check.scala 579:74:@734.4]
  wire  dat_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 579:58:@735.4]
  wire  _T_1005; // @[NV_NVDLA_CSC_dl_for_check.scala 580:39:@736.4]
  wire  _T_1006; // @[NV_NVDLA_CSC_dl_for_check.scala 580:37:@737.4]
  wire  _T_1007; // @[NV_NVDLA_CSC_dl_for_check.scala 580:56:@738.4]
  wire  dat_req_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 580:54:@739.4]
  wire  _T_1008; // @[NV_NVDLA_CSC_dl_for_check.scala 583:37:@740.4]
  wire  _T_1009; // @[NV_NVDLA_CSC_dl_for_check.scala 583:27:@741.4]
  wire  _T_1010; // @[NV_NVDLA_CSC_dl_for_check.scala 583:54:@742.4]
  wire  dat_req_sub_c_w; // @[NV_NVDLA_CSC_dl_for_check.scala 583:26:@743.4]
  wire  _T_1011; // @[NV_NVDLA_CSC_dl_for_check.scala 584:41:@744.4]
  wire  _T_1013; // @[NV_NVDLA_CSC_dl_for_check.scala 584:46:@746.4]
  wire [1:0] _T_1014; // @[NV_NVDLA_CSC_dl_for_check.scala 584:76:@747.4]
  wire [1:0] dat_req_sub_w_w; // @[NV_NVDLA_CSC_dl_for_check.scala 584:26:@748.4]
  wire  _T_1016; // @[NV_NVDLA_CSC_dl_for_check.scala 585:55:@749.4]
  wire  dat_req_sub_w_st_en; // @[NV_NVDLA_CSC_dl_for_check.scala 585:42:@750.4]
  wire  dat_req_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 588:42:@752.4]
  wire [8:0] dat_req_flag_w; // @[Cat.scala 30:58:@756.4]
  reg  dat_req_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 595:31:@757.4]
  reg [31:0] _RAND_94;
  reg [1:0] dat_req_sub_w_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 596:31:@758.4]
  reg [31:0] _RAND_95;
  reg [1:0] dat_req_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 597:31:@759.4]
  reg [31:0] _RAND_96;
  reg  dat_req_sub_c_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 598:31:@760.4]
  reg [31:0] _RAND_97;
  reg  dat_req_ch_end_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 599:32:@761.4]
  reg [31:0] _RAND_98;
  reg  dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 600:31:@762.4]
  reg [31:0] _RAND_99;
  reg [1:0] dat_req_cur_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 601:35:@763.4]
  reg [31:0] _RAND_100;
  reg  dat_req_sub_w_st_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 602:34:@764.4]
  reg [31:0] _RAND_101;
  reg [8:0] dat_req_flag_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 603:30:@765.4]
  reg [31:0] _RAND_102;
  reg  dat_req_rls_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 604:29:@766.4]
  reg [31:0] _RAND_103;
  wire  _T_1040; // @[NV_NVDLA_CSC_dl_for_check.scala 615:38:@776.6]
  wire  _T_1041; // @[NV_NVDLA_CSC_dl_for_check.scala 615:56:@777.6]
  wire [1:0] _GEN_82; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire [1:0] _GEN_83; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_84; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_85; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_86; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire [1:0] _GEN_87; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire [8:0] _GEN_88; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_89; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_90; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_91; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  wire  _GEN_92; // @[NV_NVDLA_CSC_dl_for_check.scala 619:26:@782.4]
  reg [12:0] c_bias; // @[NV_NVDLA_CSC_dl_for_check.scala 627:21:@785.4]
  reg [31:0] _RAND_104;
  reg [12:0] c_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 628:24:@786.4]
  reg [31:0] _RAND_105;
  reg [12:0] h_bias_0_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 629:26:@787.4]
  reg [31:0] _RAND_106;
  reg [12:0] h_bias_1_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 630:26:@788.4]
  reg [31:0] _RAND_107;
  reg [12:0] h_bias_2_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 631:26:@789.4]
  reg [31:0] _RAND_108;
  reg [12:0] h_bias_3_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 632:26:@790.4]
  reg [31:0] _RAND_109;
  reg [12:0] w_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 633:24:@791.4]
  reg [31:0] _RAND_110;
  wire  _T_1056; // @[NV_NVDLA_CSC_dl_for_check.scala 636:32:@792.4]
  wire  _T_1057; // @[NV_NVDLA_CSC_dl_for_check.scala 636:22:@793.4]
  wire [11:0] _T_1058; // @[NV_NVDLA_CSC_dl_for_check.scala 636:49:@794.4]
  wire [11:0] c_bias_add; // @[NV_NVDLA_CSC_dl_for_check.scala 636:21:@795.4]
  wire  _T_1061; // @[NV_NVDLA_CSC_dl_for_check.scala 638:34:@796.4]
  wire [12:0] _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 638:64:@797.4]
  wire [13:0] _T_1063; // @[NV_NVDLA_CSC_dl_for_check.scala 638:64:@797.4]
  wire [12:0] _T_1064; // @[NV_NVDLA_CSC_dl_for_check.scala 638:64:@798.4]
  wire [12:0] _T_1065; // @[NV_NVDLA_CSC_dl_for_check.scala 638:19:@799.4]
  wire [12:0] c_bias_w; // @[NV_NVDLA_CSC_dl_for_check.scala 637:19:@800.4]
  wire  c_bias_d1_reg_en; // @[NV_NVDLA_CSC_dl_for_check.scala 640:31:@804.4]
  wire [22:0] _GEN_709; // @[NV_NVDLA_CSC_dl_for_check.scala 643:32:@805.4]
  wire [36:0] _T_1068; // @[NV_NVDLA_CSC_dl_for_check.scala 643:32:@805.4]
  wire [12:0] h_bias_0_w; // @[NV_NVDLA_CSC_dl_for_check.scala 643:50:@806.4]
  wire [30:0] _GEN_710; // @[NV_NVDLA_CSC_dl_for_check.scala 644:31:@807.4]
  wire [35:0] _T_1069; // @[NV_NVDLA_CSC_dl_for_check.scala 644:31:@807.4]
  wire [12:0] h_bias_1_w; // @[NV_NVDLA_CSC_dl_for_check.scala 644:49:@808.4]
  wire [16:0] _GEN_711; // @[NV_NVDLA_CSC_dl_for_check.scala 645:29:@809.4]
  wire [21:0] _T_1070; // @[NV_NVDLA_CSC_dl_for_check.scala 645:29:@809.4]
  wire [12:0] h_bias_2_w; // @[NV_NVDLA_CSC_dl_for_check.scala 645:47:@810.4]
  wire [16:0] _GEN_712; // @[NV_NVDLA_CSC_dl_for_check.scala 646:47:@811.4]
  wire [18:0] _T_1072; // @[NV_NVDLA_CSC_dl_for_check.scala 646:47:@811.4]
  wire [18:0] _T_1073; // @[NV_NVDLA_CSC_dl_for_check.scala 646:21:@812.4]
  wire [12:0] h_bias_3_w; // @[NV_NVDLA_CSC_dl_for_check.scala 646:65:@813.4]
  wire  _T_1074; // @[NV_NVDLA_CSC_dl_for_check.scala 647:69:@814.4]
  wire  _T_1075; // @[NV_NVDLA_CSC_dl_for_check.scala 647:84:@815.4]
  wire  _T_1076; // @[NV_NVDLA_CSC_dl_for_check.scala 647:73:@816.4]
  wire  _T_1077; // @[NV_NVDLA_CSC_dl_for_check.scala 647:52:@817.4]
  wire  _T_1078; // @[NV_NVDLA_CSC_dl_for_check.scala 647:34:@818.4]
  wire [1:0] h_bias_reg_en; // @[Cat.scala 30:58:@819.4]
  wire [12:0] _GEN_93; // @[NV_NVDLA_CSC_dl_for_check.scala 677:20:@840.4]
  wire [12:0] _GEN_94; // @[NV_NVDLA_CSC_dl_for_check.scala 680:23:@843.4]
  wire  _T_1101; // @[NV_NVDLA_CSC_dl_for_check.scala 683:19:@846.4]
  wire [12:0] _GEN_95; // @[NV_NVDLA_CSC_dl_for_check.scala 683:23:@847.4]
  wire [12:0] _GEN_96; // @[NV_NVDLA_CSC_dl_for_check.scala 683:23:@847.4]
  wire [12:0] _GEN_97; // @[NV_NVDLA_CSC_dl_for_check.scala 683:23:@847.4]
  wire  _T_1102; // @[NV_NVDLA_CSC_dl_for_check.scala 688:19:@852.4]
  wire [12:0] _GEN_98; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@853.4]
  wire [13:0] _GEN_99; // @[NV_NVDLA_CSC_dl_for_check.scala 691:20:@856.4]
  reg [12:0] dat_req_sub_h_addr_0; // @[NV_NVDLA_CSC_dl_for_check.scala 699:33:@868.4]
  reg [31:0] _RAND_111;
  reg [12:0] dat_req_sub_h_addr_1; // @[NV_NVDLA_CSC_dl_for_check.scala 699:33:@868.4]
  reg [31:0] _RAND_112;
  reg [12:0] dat_req_sub_h_addr_2; // @[NV_NVDLA_CSC_dl_for_check.scala 699:33:@868.4]
  reg [31:0] _RAND_113;
  reg [12:0] dat_req_sub_h_addr_3; // @[NV_NVDLA_CSC_dl_for_check.scala 699:33:@868.4]
  reg [31:0] _RAND_114;
  reg  sc2buf_dat_rd_en_out; // @[NV_NVDLA_CSC_dl_for_check.scala 700:35:@869.4]
  reg [31:0] _RAND_115;
  reg [18:0] sc2buf_dat_rd_addr_out; // @[NV_NVDLA_CSC_dl_for_check.scala 701:37:@871.4]
  reg [31:0] _RAND_116;
  reg  dat_req_pipe_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 702:32:@872.4]
  reg [31:0] _RAND_117;
  reg  dat_req_exec_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 703:32:@873.4]
  reg [31:0] _RAND_118;
  reg  dat_req_exec_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 705:33:@875.4]
  reg [31:0] _RAND_119;
  reg [1:0] dat_req_pipe_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 706:33:@876.4]
  reg [31:0] _RAND_120;
  reg [1:0] dat_req_pipe_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 707:33:@877.4]
  reg [31:0] _RAND_121;
  reg  dat_req_pipe_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 708:33:@878.4]
  reg [31:0] _RAND_122;
  reg  dat_req_pipe_ch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 709:34:@879.4]
  reg [31:0] _RAND_123;
  reg [7:0] dat_req_pipe_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 710:33:@880.4]
  reg [31:0] _RAND_124;
  reg  dat_req_pipe_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 711:33:@881.4]
  reg [31:0] _RAND_125;
  reg [1:0] dat_req_pipe_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 712:37:@882.4]
  reg [31:0] _RAND_126;
  reg  dat_req_pipe_sub_w_st; // @[NV_NVDLA_CSC_dl_for_check.scala 713:36:@883.4]
  reg [31:0] _RAND_127;
  reg  dat_req_pipe_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 714:31:@884.4]
  reg [31:0] _RAND_128;
  reg [8:0] dat_req_pipe_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 715:32:@885.4]
  reg [31:0] _RAND_129;
  wire [13:0] _T_1197; // @[NV_NVDLA_CSC_dl_for_check.scala 717:30:@886.4]
  wire [13:0] _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 717:45:@887.4]
  wire [14:0] _T_1198; // @[NV_NVDLA_CSC_dl_for_check.scala 717:45:@887.4]
  wire [14:0] _GEN_714; // @[NV_NVDLA_CSC_dl_for_check.scala 717:60:@888.4]
  wire [15:0] _T_1199; // @[NV_NVDLA_CSC_dl_for_check.scala 717:60:@888.4]
  wire [12:0] h_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 717:75:@889.4]
  wire [14:0] _GEN_715; // @[NV_NVDLA_CSC_dl_for_check.scala 718:40:@890.4]
  wire [15:0] _T_1200; // @[NV_NVDLA_CSC_dl_for_check.scala 718:40:@890.4]
  wire [15:0] _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 718:53:@891.4]
  wire [16:0] _T_1201; // @[NV_NVDLA_CSC_dl_for_check.scala 718:53:@891.4]
  wire [16:0] _GEN_717; // @[NV_NVDLA_CSC_dl_for_check.scala 718:66:@892.4]
  wire [17:0] dat_req_addr_sum; // @[NV_NVDLA_CSC_dl_for_check.scala 718:66:@892.4]
  wire [17:0] _GEN_718; // @[NV_NVDLA_CSC_dl_for_check.scala 719:45:@895.4]
  wire  is_dat_req_addr_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 719:45:@895.4]
  wire [18:0] _T_1214; // @[NV_NVDLA_CSC_dl_for_check.scala 720:42:@898.4]
  wire [18:0] dat_req_addr_wrap; // @[NV_NVDLA_CSC_dl_for_check.scala 720:42:@899.4]
  wire  _T_1215; // @[NV_NVDLA_CSC_dl_for_check.scala 721:35:@900.4]
  wire [18:0] _T_1221; // @[NV_NVDLA_CSC_dl_for_check.scala 722:25:@902.4]
  wire [18:0] dat_req_addr_w; // @[NV_NVDLA_CSC_dl_for_check.scala 721:25:@903.4]
  wire  _T_1225; // @[Mux.scala 46:19:@904.4]
  wire [12:0] _T_1226; // @[Mux.scala 46:16:@905.4]
  wire  _T_1227; // @[Mux.scala 46:19:@906.4]
  wire [12:0] _T_1228; // @[Mux.scala 46:16:@907.4]
  wire  _T_1229; // @[Mux.scala 46:19:@908.4]
  wire [12:0] dat_req_addr_last; // @[Mux.scala 46:16:@909.4]
  wire [18:0] _GEN_720; // @[NV_NVDLA_CSC_dl_for_check.scala 725:65:@910.4]
  wire  _T_1230; // @[NV_NVDLA_CSC_dl_for_check.scala 725:65:@910.4]
  wire  _T_1231; // @[NV_NVDLA_CSC_dl_for_check.scala 725:85:@911.4]
  wire  sc2buf_dat_rd_en_w; // @[NV_NVDLA_CSC_dl_for_check.scala 725:43:@912.4]
  wire  _T_1232; // @[NV_NVDLA_CSC_dl_for_check.scala 727:38:@913.4]
  wire  _T_1234; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@914.4]
  wire  _T_1235; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@915.4]
  wire  dat_req_sub_h_addr_en_0; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@916.4]
  wire  _T_1239; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@918.4]
  wire  _T_1240; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@919.4]
  wire  dat_req_sub_h_addr_en_1; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@920.4]
  wire  _T_1244; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@922.4]
  wire  _T_1245; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@923.4]
  wire  dat_req_sub_h_addr_en_2; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@924.4]
  wire  _T_1249; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@926.4]
  wire  _T_1250; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@927.4]
  wire  dat_req_sub_h_addr_en_3; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@928.4]
  wire [18:0] _GEN_100; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@934.4]
  wire [18:0] _GEN_101; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@937.4]
  wire [18:0] _GEN_102; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@940.4]
  wire [18:0] _GEN_103; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@943.4]
  wire  _T_1261; // @[NV_NVDLA_CSC_dl_for_check.scala 740:14:@947.4]
  wire [18:0] _GEN_104; // @[NV_NVDLA_CSC_dl_for_check.scala 740:34:@948.4]
  wire [1:0] _GEN_105; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire [1:0] _GEN_106; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire  _GEN_107; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire  _GEN_108; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire [7:0] _GEN_109; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire  _GEN_110; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire [1:0] _GEN_111; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire  _GEN_112; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire  _GEN_113; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire [8:0] _GEN_114; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire  _GEN_115; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  wire [6:0] _T_1266; // @[Cat.scala 30:58:@971.4]
  wire [28:0] dat_req_pipe_pd; // @[Cat.scala 30:58:@977.4]
  reg  _T_1276; // @[NV_NVDLA_CSC_dl_for_check.scala 774:73:@979.4]
  reg [31:0] _RAND_130;
  reg  _T_1279; // @[NV_NVDLA_CSC_dl_for_check.scala 774:73:@980.4]
  reg [31:0] _RAND_131;
  reg  _T_1282; // @[NV_NVDLA_CSC_dl_for_check.scala 774:73:@981.4]
  reg [31:0] _RAND_132;
  reg  _T_1285; // @[NV_NVDLA_CSC_dl_for_check.scala 774:73:@982.4]
  reg [31:0] _RAND_133;
  reg  _T_1288; // @[NV_NVDLA_CSC_dl_for_check.scala 774:73:@983.4]
  reg [31:0] _RAND_134;
  reg  dat_rsp_pipe_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 774:73:@984.4]
  reg [31:0] _RAND_135;
  reg [28:0] _T_1295; // @[NV_NVDLA_CSC_dl_for_check.scala 776:71:@986.4]
  reg [31:0] _RAND_136;
  reg [28:0] _T_1298; // @[NV_NVDLA_CSC_dl_for_check.scala 776:71:@987.4]
  reg [31:0] _RAND_137;
  reg [28:0] _T_1301; // @[NV_NVDLA_CSC_dl_for_check.scala 776:71:@988.4]
  reg [31:0] _RAND_138;
  reg [28:0] _T_1304; // @[NV_NVDLA_CSC_dl_for_check.scala 776:71:@989.4]
  reg [31:0] _RAND_139;
  reg [28:0] _T_1307; // @[NV_NVDLA_CSC_dl_for_check.scala 776:71:@990.4]
  reg [31:0] _RAND_140;
  reg [28:0] dat_rsp_pipe_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 776:71:@991.4]
  reg [31:0] _RAND_141;
  reg  _T_1314; // @[NV_NVDLA_CSC_dl_for_check.scala 778:73:@993.4]
  reg [31:0] _RAND_142;
  reg  _T_1317; // @[NV_NVDLA_CSC_dl_for_check.scala 778:73:@994.4]
  reg [31:0] _RAND_143;
  reg  _T_1320; // @[NV_NVDLA_CSC_dl_for_check.scala 778:73:@995.4]
  reg [31:0] _RAND_144;
  reg  _T_1323; // @[NV_NVDLA_CSC_dl_for_check.scala 778:73:@996.4]
  reg [31:0] _RAND_145;
  reg  _T_1326; // @[NV_NVDLA_CSC_dl_for_check.scala 778:73:@997.4]
  reg [31:0] _RAND_146;
  reg  dat_rsp_exec_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 778:73:@998.4]
  reg [31:0] _RAND_147;
  reg  _T_1333; // @[NV_NVDLA_CSC_dl_for_check.scala 780:73:@1000.4]
  reg [31:0] _RAND_148;
  reg  _T_1336; // @[NV_NVDLA_CSC_dl_for_check.scala 780:73:@1001.4]
  reg [31:0] _RAND_149;
  reg  _T_1339; // @[NV_NVDLA_CSC_dl_for_check.scala 780:73:@1002.4]
  reg [31:0] _RAND_150;
  reg  _T_1342; // @[NV_NVDLA_CSC_dl_for_check.scala 780:73:@1003.4]
  reg [31:0] _RAND_151;
  reg  _T_1345; // @[NV_NVDLA_CSC_dl_for_check.scala 780:73:@1004.4]
  reg [31:0] _RAND_152;
  reg  dat_rsp_exec_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 780:73:@1005.4]
  reg [31:0] _RAND_153;
  reg [1:0] _T_1352; // @[NV_NVDLA_CSC_dl_for_check.scala 782:74:@1007.4]
  reg [31:0] _RAND_154;
  reg [1:0] _T_1355; // @[NV_NVDLA_CSC_dl_for_check.scala 782:74:@1008.4]
  reg [31:0] _RAND_155;
  reg [1:0] _T_1358; // @[NV_NVDLA_CSC_dl_for_check.scala 782:74:@1009.4]
  reg [31:0] _RAND_156;
  reg [1:0] _T_1361; // @[NV_NVDLA_CSC_dl_for_check.scala 782:74:@1010.4]
  reg [31:0] _RAND_157;
  reg [1:0] _T_1364; // @[NV_NVDLA_CSC_dl_for_check.scala 782:74:@1011.4]
  reg [31:0] _RAND_158;
  reg [1:0] dat_rsp_exec_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 782:74:@1012.4]
  reg [31:0] _RAND_159;
  wire [28:0] _GEN_116; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1019.4]
  wire  _GEN_117; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1023.4]
  wire [1:0] _GEN_118; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1023.4]
  wire [28:0] _GEN_119; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1028.4]
  wire  _GEN_120; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1032.4]
  wire [1:0] _GEN_121; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1032.4]
  wire [28:0] _GEN_122; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1037.4]
  wire  _GEN_123; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1041.4]
  wire [1:0] _GEN_124; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1041.4]
  wire [28:0] _GEN_125; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1046.4]
  wire  _GEN_126; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1050.4]
  wire [1:0] _GEN_127; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1050.4]
  wire [28:0] _GEN_128; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1055.4]
  wire  _GEN_129; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1059.4]
  wire [1:0] _GEN_130; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1059.4]
  wire [28:0] _GEN_131; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1064.4]
  wire  _GEN_132; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1068.4]
  wire [1:0] _GEN_133; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1068.4]
  wire [1:0] dat_rsp_pipe_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 809:41:@1072.4]
  wire [1:0] dat_rsp_pipe_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 810:41:@1073.4]
  wire  dat_rsp_pipe_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 811:41:@1074.4]
  wire  dat_rsp_pipe_ch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 812:42:@1075.4]
  wire [7:0] dat_rsp_pipe_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 813:41:@1076.4]
  wire [1:0] dat_rsp_pipe_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 814:45:@1077.4]
  wire  dat_rsp_pipe_sub_w_st; // @[NV_NVDLA_CSC_dl_for_check.scala 816:44:@1079.4]
  wire  dat_rsp_pipe_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 817:39:@1080.4]
  wire [8:0] dat_rsp_pipe_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 818:40:@1081.4]
  reg  dat_l0c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 823:29:@1082.4]
  reg [31:0] _RAND_160;
  reg  dat_l1c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 824:29:@1083.4]
  reg [31:0] _RAND_161;
  reg  dat_l2c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 825:29:@1084.4]
  reg [31:0] _RAND_162;
  reg  dat_l3c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 826:29:@1085.4]
  reg [31:0] _RAND_163;
  reg  dat_l0c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 827:29:@1086.4]
  reg [31:0] _RAND_164;
  reg  dat_l1c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 828:29:@1087.4]
  reg [31:0] _RAND_165;
  reg  dat_l2c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 829:29:@1088.4]
  reg [31:0] _RAND_166;
  reg  dat_l3c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 830:29:@1089.4]
  reg [31:0] _RAND_167;
  reg [511:0] dat_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 832:19:@1090.4]
  reg [511:0] _RAND_168;
  reg [511:0] dat_l1c0; // @[NV_NVDLA_CSC_dl_for_check.scala 833:19:@1091.4]
  reg [511:0] _RAND_169;
  reg [511:0] dat_l2c0; // @[NV_NVDLA_CSC_dl_for_check.scala 834:19:@1092.4]
  reg [511:0] _RAND_170;
  reg [511:0] dat_l3c0; // @[NV_NVDLA_CSC_dl_for_check.scala 835:19:@1093.4]
  reg [511:0] _RAND_171;
  reg [511:0] dat_l0c1; // @[NV_NVDLA_CSC_dl_for_check.scala 836:19:@1094.4]
  reg [511:0] _RAND_172;
  reg [511:0] dat_l1c1; // @[NV_NVDLA_CSC_dl_for_check.scala 837:19:@1095.4]
  reg [511:0] _RAND_173;
  reg [511:0] dat_l2c1; // @[NV_NVDLA_CSC_dl_for_check.scala 838:19:@1096.4]
  reg [511:0] _RAND_174;
  reg [511:0] dat_l3c1; // @[NV_NVDLA_CSC_dl_for_check.scala 839:19:@1097.4]
  reg [511:0] _RAND_175;
  wire  _T_1392; // @[NV_NVDLA_CSC_dl_for_check.scala 841:70:@1098.4]
  wire  dat_l0c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 841:48:@1099.4]
  wire  _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 842:70:@1100.4]
  wire  dat_l1c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 842:48:@1101.4]
  wire  _T_1396; // @[NV_NVDLA_CSC_dl_for_check.scala 843:70:@1102.4]
  wire  dat_l2c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 843:48:@1103.4]
  wire  _T_1398; // @[NV_NVDLA_CSC_dl_for_check.scala 844:70:@1104.4]
  wire  dat_l3c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 844:48:@1105.4]
  wire  _T_1399; // @[NV_NVDLA_CSC_dl_for_check.scala 847:62:@1106.4]
  wire  _T_1400; // @[NV_NVDLA_CSC_dl_for_check.scala 847:46:@1107.4]
  wire  _T_1401; // @[NV_NVDLA_CSC_dl_for_check.scala 847:69:@1108.4]
  wire  dat_wg_adv; // @[NV_NVDLA_CSC_dl_for_check.scala 847:67:@1109.4]
  wire  _T_1402; // @[NV_NVDLA_CSC_dl_for_check.scala 848:52:@1110.4]
  wire  _T_1403; // @[NV_NVDLA_CSC_dl_for_check.scala 848:33:@1111.4]
  wire  _T_1404; // @[NV_NVDLA_CSC_dl_for_check.scala 848:31:@1112.4]
  wire  _T_1405; // @[NV_NVDLA_CSC_dl_for_check.scala 848:69:@1113.4]
  wire  _T_1406; // @[NV_NVDLA_CSC_dl_for_check.scala 848:74:@1114.4]
  wire  _T_1407; // @[NV_NVDLA_CSC_dl_for_check.scala 848:90:@1115.4]
  wire  _T_1408; // @[NV_NVDLA_CSC_dl_for_check.scala 848:88:@1116.4]
  wire  dat_l0c1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 848:57:@1117.4]
  wire  _T_1410; // @[NV_NVDLA_CSC_dl_for_check.scala 849:31:@1119.4]
  wire  _T_1411; // @[NV_NVDLA_CSC_dl_for_check.scala 849:68:@1120.4]
  wire  _T_1412; // @[NV_NVDLA_CSC_dl_for_check.scala 849:73:@1121.4]
  wire  _T_1413; // @[NV_NVDLA_CSC_dl_for_check.scala 849:89:@1122.4]
  wire  _T_1414; // @[NV_NVDLA_CSC_dl_for_check.scala 849:87:@1123.4]
  wire  dat_l1c1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 849:56:@1124.4]
  wire  _T_1415; // @[NV_NVDLA_CSC_dl_for_check.scala 850:29:@1125.4]
  wire  _T_1416; // @[NV_NVDLA_CSC_dl_for_check.scala 850:34:@1126.4]
  wire  _T_1417; // @[NV_NVDLA_CSC_dl_for_check.scala 850:50:@1127.4]
  wire  dat_l2c1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 850:48:@1128.4]
  wire  _T_1418; // @[NV_NVDLA_CSC_dl_for_check.scala 851:29:@1129.4]
  wire  _T_1419; // @[NV_NVDLA_CSC_dl_for_check.scala 851:34:@1130.4]
  wire  _T_1420; // @[NV_NVDLA_CSC_dl_for_check.scala 851:50:@1131.4]
  wire  dat_l3c1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 851:48:@1132.4]
  wire  _T_1421; // @[NV_NVDLA_CSC_dl_for_check.scala 853:41:@1133.4]
  wire  dat_dummy_l0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 853:62:@1135.4]
  wire  dat_dummy_l1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 854:62:@1138.4]
  wire  dat_dummy_l2_en; // @[NV_NVDLA_CSC_dl_for_check.scala 855:62:@1141.4]
  wire  dat_dummy_l3_en; // @[NV_NVDLA_CSC_dl_for_check.scala 856:62:@1144.4]
  wire  dat_l0_set; // @[NV_NVDLA_CSC_dl_for_check.scala 858:30:@1145.4]
  wire  dat_l1_set; // @[NV_NVDLA_CSC_dl_for_check.scala 859:30:@1146.4]
  wire  dat_l2_set; // @[NV_NVDLA_CSC_dl_for_check.scala 860:30:@1147.4]
  wire  dat_l3_set; // @[NV_NVDLA_CSC_dl_for_check.scala 861:30:@1148.4]
  wire  _T_1435; // @[NV_NVDLA_CSC_dl_for_check.scala 863:48:@1149.4]
  wire  _T_1436; // @[NV_NVDLA_CSC_dl_for_check.scala 863:22:@1150.4]
  wire  _T_1439; // @[NV_NVDLA_CSC_dl_for_check.scala 864:48:@1152.4]
  wire  _T_1440; // @[NV_NVDLA_CSC_dl_for_check.scala 864:22:@1153.4]
  wire  _T_1443; // @[NV_NVDLA_CSC_dl_for_check.scala 865:48:@1155.4]
  wire  _T_1444; // @[NV_NVDLA_CSC_dl_for_check.scala 865:22:@1156.4]
  wire  _T_1447; // @[NV_NVDLA_CSC_dl_for_check.scala 866:48:@1158.4]
  wire  _T_1448; // @[NV_NVDLA_CSC_dl_for_check.scala 866:22:@1159.4]
  wire  _T_1450; // @[NV_NVDLA_CSC_dl_for_check.scala 867:48:@1161.4]
  wire  _T_1451; // @[NV_NVDLA_CSC_dl_for_check.scala 867:22:@1162.4]
  wire  _T_1454; // @[NV_NVDLA_CSC_dl_for_check.scala 868:77:@1164.4]
  wire  _T_1455; // @[NV_NVDLA_CSC_dl_for_check.scala 868:60:@1165.4]
  wire  _T_1456; // @[NV_NVDLA_CSC_dl_for_check.scala 868:48:@1166.4]
  wire  _T_1457; // @[NV_NVDLA_CSC_dl_for_check.scala 868:22:@1167.4]
  wire  _T_1459; // @[NV_NVDLA_CSC_dl_for_check.scala 869:76:@1169.4]
  wire  _T_1460; // @[NV_NVDLA_CSC_dl_for_check.scala 869:60:@1170.4]
  wire  _T_1461; // @[NV_NVDLA_CSC_dl_for_check.scala 869:48:@1171.4]
  wire  _T_1462; // @[NV_NVDLA_CSC_dl_for_check.scala 869:22:@1172.4]
  wire  _T_1465; // @[NV_NVDLA_CSC_dl_for_check.scala 870:60:@1175.4]
  wire  _T_1466; // @[NV_NVDLA_CSC_dl_for_check.scala 870:48:@1176.4]
  wire  _T_1467; // @[NV_NVDLA_CSC_dl_for_check.scala 870:22:@1177.4]
  reg [7:0] rsp_sft_cnt_l0; // @[NV_NVDLA_CSC_dl_for_check.scala 884:29:@1203.4]
  reg [31:0] _RAND_176;
  reg [7:0] rsp_sft_cnt_l1; // @[NV_NVDLA_CSC_dl_for_check.scala 885:29:@1204.4]
  reg [31:0] _RAND_177;
  reg [7:0] rsp_sft_cnt_l2; // @[NV_NVDLA_CSC_dl_for_check.scala 886:29:@1205.4]
  reg [31:0] _RAND_178;
  reg [7:0] rsp_sft_cnt_l3; // @[NV_NVDLA_CSC_dl_for_check.scala 887:29:@1206.4]
  reg [31:0] _RAND_179;
  reg [7:0] rsp_sft_cnt_l0_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 888:33:@1207.4]
  reg [31:0] _RAND_180;
  reg [7:0] rsp_sft_cnt_l1_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 889:33:@1208.4]
  reg [31:0] _RAND_181;
  reg [7:0] rsp_sft_cnt_l2_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 890:33:@1209.4]
  reg [31:0] _RAND_182;
  reg [7:0] rsp_sft_cnt_l3_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 891:33:@1210.4]
  reg [31:0] _RAND_183;
  reg  dat_rsp_l2_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 896:41:@1214.4]
  reg [31:0] _RAND_184;
  reg [26:0] _T_1504; // @[NV_NVDLA_CSC_dl_for_check.scala 898:41:@1219.4]
  reg [31:0] _RAND_185;
  wire [26:0] _T_1516; // @[Cat.scala 30:58:@1229.4]
  wire [26:0] _GEN_142; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1232.4]
  wire [26:0] _GEN_143; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1236.4]
  wire [26:0] _GEN_144; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1240.4]
  wire [26:0] _GEN_145; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1244.4]
  wire  dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 924:39:@1270.4]
  wire  dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 925:39:@1271.4]
  wire  dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 926:39:@1272.4]
  wire  dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 927:39:@1273.4]
  wire [8:0] dat_rsp_l0_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 929:38:@1274.4]
  wire [8:0] dat_rsp_l1_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 930:38:@1275.4]
  wire [8:0] dat_rsp_l2_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 931:38:@1276.4]
  wire [8:0] dat_rsp_l3_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 932:38:@1277.4]
  wire  dat_rsp_l0_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 934:44:@1278.4]
  wire  dat_rsp_l1_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 935:44:@1279.4]
  wire  dat_rsp_l2_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 936:44:@1280.4]
  wire  dat_rsp_l3_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 937:44:@1281.4]
  wire [1:0] dat_rsp_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 940:31:@1282.4]
  wire [7:0] dat_rsp_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 944:31:@1286.4]
  wire [1:0] dat_rsp_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 945:35:@1287.4]
  wire [8:0] dat_rsp_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 947:30:@1290.4]
  wire [7:0] rsp_sft_cnt_l0_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 956:29:@1296.4]
  wire [7:0] rsp_sft_cnt_l1_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 957:29:@1297.4]
  wire [7:0] rsp_sft_cnt_l2_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 958:29:@1298.4]
  wire [7:0] rsp_sft_cnt_l3_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 959:29:@1299.4]
  wire  _T_1554; // @[NV_NVDLA_CSC_dl_for_check.scala 961:50:@1300.4]
  wire [7:0] _GEN_721; // @[NV_NVDLA_CSC_dl_for_check.scala 961:111:@1301.4]
  wire [8:0] _T_1556; // @[NV_NVDLA_CSC_dl_for_check.scala 961:111:@1301.4]
  wire [8:0] _GEN_722; // @[NV_NVDLA_CSC_dl_for_check.scala 961:134:@1302.4]
  wire [9:0] _T_1557; // @[NV_NVDLA_CSC_dl_for_check.scala 961:134:@1302.4]
  wire [9:0] _T_1558; // @[NV_NVDLA_CSC_dl_for_check.scala 961:134:@1303.4]
  wire [9:0] _T_1559; // @[NV_NVDLA_CSC_dl_for_check.scala 961:29:@1304.4]
  wire [7:0] rsp_sft_cnt_l0_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 961:156:@1305.4]
  wire [8:0] _T_1563; // @[NV_NVDLA_CSC_dl_for_check.scala 962:111:@1307.4]
  wire [8:0] _GEN_724; // @[NV_NVDLA_CSC_dl_for_check.scala 962:134:@1308.4]
  wire [9:0] _T_1564; // @[NV_NVDLA_CSC_dl_for_check.scala 962:134:@1308.4]
  wire [9:0] _T_1565; // @[NV_NVDLA_CSC_dl_for_check.scala 962:134:@1309.4]
  wire [9:0] _T_1566; // @[NV_NVDLA_CSC_dl_for_check.scala 962:29:@1310.4]
  wire [7:0] rsp_sft_cnt_l1_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 962:156:@1311.4]
  wire [8:0] _T_1570; // @[NV_NVDLA_CSC_dl_for_check.scala 963:111:@1313.4]
  wire [8:0] _GEN_726; // @[NV_NVDLA_CSC_dl_for_check.scala 963:134:@1314.4]
  wire [9:0] _T_1571; // @[NV_NVDLA_CSC_dl_for_check.scala 963:134:@1314.4]
  wire [9:0] _T_1572; // @[NV_NVDLA_CSC_dl_for_check.scala 963:134:@1315.4]
  wire [9:0] _T_1573; // @[NV_NVDLA_CSC_dl_for_check.scala 963:29:@1316.4]
  wire [7:0] rsp_sft_cnt_l2_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 963:156:@1317.4]
  wire [8:0] _T_1577; // @[NV_NVDLA_CSC_dl_for_check.scala 964:111:@1319.4]
  wire [8:0] _GEN_728; // @[NV_NVDLA_CSC_dl_for_check.scala 964:134:@1320.4]
  wire [9:0] _T_1578; // @[NV_NVDLA_CSC_dl_for_check.scala 964:134:@1320.4]
  wire [9:0] _T_1579; // @[NV_NVDLA_CSC_dl_for_check.scala 964:134:@1321.4]
  wire [9:0] _T_1580; // @[NV_NVDLA_CSC_dl_for_check.scala 964:29:@1322.4]
  wire [7:0] rsp_sft_cnt_l3_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 964:156:@1323.4]
  wire  _T_1582; // @[NV_NVDLA_CSC_dl_for_check.scala 973:52:@1324.4]
  wire  _T_1583; // @[NV_NVDLA_CSC_dl_for_check.scala 973:50:@1325.4]
  wire  _T_1584; // @[NV_NVDLA_CSC_dl_for_check.scala 974:50:@1326.4]
  wire [7:0] _T_1587; // @[NV_NVDLA_CSC_dl_for_check.scala 975:64:@1327.4]
  wire [7:0] _T_1588; // @[NV_NVDLA_CSC_dl_for_check.scala 975:27:@1328.4]
  wire [7:0] _T_1589; // @[NV_NVDLA_CSC_dl_for_check.scala 974:27:@1329.4]
  wire [7:0] _T_1590; // @[NV_NVDLA_CSC_dl_for_check.scala 973:27:@1330.4]
  wire [7:0] rsp_sft_cnt_l0_w; // @[NV_NVDLA_CSC_dl_for_check.scala 972:27:@1331.4]
  wire  _T_1592; // @[NV_NVDLA_CSC_dl_for_check.scala 978:52:@1332.4]
  wire  _T_1593; // @[NV_NVDLA_CSC_dl_for_check.scala 978:50:@1333.4]
  wire  _T_1594; // @[NV_NVDLA_CSC_dl_for_check.scala 979:50:@1334.4]
  wire [7:0] _T_1597; // @[NV_NVDLA_CSC_dl_for_check.scala 980:64:@1335.4]
  wire [7:0] _T_1598; // @[NV_NVDLA_CSC_dl_for_check.scala 980:27:@1336.4]
  wire [7:0] _T_1599; // @[NV_NVDLA_CSC_dl_for_check.scala 979:27:@1337.4]
  wire [7:0] _T_1600; // @[NV_NVDLA_CSC_dl_for_check.scala 978:27:@1338.4]
  wire [7:0] rsp_sft_cnt_l1_w; // @[NV_NVDLA_CSC_dl_for_check.scala 977:27:@1339.4]
  wire  _T_1602; // @[NV_NVDLA_CSC_dl_for_check.scala 983:52:@1340.4]
  wire  _T_1603; // @[NV_NVDLA_CSC_dl_for_check.scala 983:50:@1341.4]
  wire  _T_1604; // @[NV_NVDLA_CSC_dl_for_check.scala 984:50:@1342.4]
  wire [7:0] _T_1607; // @[NV_NVDLA_CSC_dl_for_check.scala 985:64:@1343.4]
  wire [7:0] _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 985:27:@1344.4]
  wire [7:0] _T_1609; // @[NV_NVDLA_CSC_dl_for_check.scala 984:27:@1345.4]
  wire [7:0] _T_1610; // @[NV_NVDLA_CSC_dl_for_check.scala 983:27:@1346.4]
  wire [7:0] rsp_sft_cnt_l2_w; // @[NV_NVDLA_CSC_dl_for_check.scala 982:27:@1347.4]
  wire  _T_1612; // @[NV_NVDLA_CSC_dl_for_check.scala 988:52:@1348.4]
  wire  _T_1613; // @[NV_NVDLA_CSC_dl_for_check.scala 988:50:@1349.4]
  wire  _T_1614; // @[NV_NVDLA_CSC_dl_for_check.scala 989:50:@1350.4]
  wire [7:0] _T_1617; // @[NV_NVDLA_CSC_dl_for_check.scala 990:64:@1351.4]
  wire [7:0] _T_1618; // @[NV_NVDLA_CSC_dl_for_check.scala 990:27:@1352.4]
  wire [7:0] _T_1619; // @[NV_NVDLA_CSC_dl_for_check.scala 989:27:@1353.4]
  wire [7:0] _T_1620; // @[NV_NVDLA_CSC_dl_for_check.scala 988:27:@1354.4]
  wire [7:0] rsp_sft_cnt_l3_w; // @[NV_NVDLA_CSC_dl_for_check.scala 987:27:@1355.4]
  wire  _T_1621; // @[NV_NVDLA_CSC_dl_for_check.scala 993:46:@1356.4]
  wire  _T_1622; // @[NV_NVDLA_CSC_dl_for_check.scala 993:51:@1357.4]
  wire  rsp_sft_cnt_l0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 993:34:@1358.4]
  wire  _T_1623; // @[NV_NVDLA_CSC_dl_for_check.scala 994:46:@1359.4]
  wire  _T_1624; // @[NV_NVDLA_CSC_dl_for_check.scala 994:51:@1360.4]
  wire  _T_1626; // @[NV_NVDLA_CSC_dl_for_check.scala 994:87:@1361.4]
  wire  _T_1627; // @[NV_NVDLA_CSC_dl_for_check.scala 994:69:@1362.4]
  wire  rsp_sft_cnt_l1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 994:34:@1363.4]
  wire  _T_1628; // @[NV_NVDLA_CSC_dl_for_check.scala 995:46:@1364.4]
  wire  _T_1629; // @[NV_NVDLA_CSC_dl_for_check.scala 995:51:@1365.4]
  wire  _T_1631; // @[NV_NVDLA_CSC_dl_for_check.scala 995:87:@1366.4]
  wire  _T_1632; // @[NV_NVDLA_CSC_dl_for_check.scala 995:69:@1367.4]
  wire  rsp_sft_cnt_l2_en; // @[NV_NVDLA_CSC_dl_for_check.scala 995:34:@1368.4]
  wire  _T_1633; // @[NV_NVDLA_CSC_dl_for_check.scala 996:46:@1369.4]
  wire  _T_1634; // @[NV_NVDLA_CSC_dl_for_check.scala 996:51:@1370.4]
  wire  _T_1637; // @[NV_NVDLA_CSC_dl_for_check.scala 996:69:@1372.4]
  wire  rsp_sft_cnt_l3_en; // @[NV_NVDLA_CSC_dl_for_check.scala 996:34:@1373.4]
  wire  _T_1638; // @[NV_NVDLA_CSC_dl_for_check.scala 998:50:@1374.4]
  wire  _T_1639; // @[NV_NVDLA_CSC_dl_for_check.scala 998:55:@1375.4]
  wire  _T_1640; // @[NV_NVDLA_CSC_dl_for_check.scala 998:73:@1376.4]
  wire  _T_1641; // @[NV_NVDLA_CSC_dl_for_check.scala 998:97:@1377.4]
  wire  rsp_sft_cnt_l0_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 998:38:@1378.4]
  wire  _T_1642; // @[NV_NVDLA_CSC_dl_for_check.scala 999:50:@1379.4]
  wire  _T_1643; // @[NV_NVDLA_CSC_dl_for_check.scala 999:55:@1380.4]
  wire  _T_1644; // @[NV_NVDLA_CSC_dl_for_check.scala 999:73:@1381.4]
  wire  _T_1645; // @[NV_NVDLA_CSC_dl_for_check.scala 999:97:@1382.4]
  wire  _T_1647; // @[NV_NVDLA_CSC_dl_for_check.scala 999:138:@1383.4]
  wire  _T_1648; // @[NV_NVDLA_CSC_dl_for_check.scala 999:120:@1384.4]
  wire  rsp_sft_cnt_l1_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 999:38:@1385.4]
  wire  _T_1649; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:50:@1386.4]
  wire  _T_1650; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:55:@1387.4]
  wire  _T_1651; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:73:@1388.4]
  wire  _T_1652; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:97:@1389.4]
  wire  _T_1654; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:138:@1390.4]
  wire  _T_1655; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:120:@1391.4]
  wire  rsp_sft_cnt_l2_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:38:@1392.4]
  wire  _T_1656; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:50:@1393.4]
  wire  _T_1657; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:55:@1394.4]
  wire  _T_1658; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:73:@1395.4]
  wire  _T_1659; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:97:@1396.4]
  wire  _T_1662; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:120:@1398.4]
  wire  rsp_sft_cnt_l3_ori_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:38:@1399.4]
  wire [7:0] _GEN_146; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:24:@1400.4]
  wire [7:0] _GEN_147; // @[NV_NVDLA_CSC_dl_for_check.scala 1004:24:@1403.4]
  wire [7:0] _GEN_148; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:24:@1406.4]
  wire [7:0] _GEN_149; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:24:@1409.4]
  wire [7:0] _GEN_150; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:28:@1412.4]
  wire [7:0] _GEN_151; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:28:@1415.4]
  wire [7:0] _GEN_152; // @[NV_NVDLA_CSC_dl_for_check.scala 1009:28:@1418.4]
  wire [7:0] _GEN_153; // @[NV_NVDLA_CSC_dl_for_check.scala 1010:28:@1421.4]
  wire [7:0] _T_1663; // @[NV_NVDLA_CSC_dl_for_check.scala 1019:55:@1424.4]
  wire [63:0] _T_1666; // @[Cat.scala 30:58:@1427.4]
  wire [127:0] _T_1667; // @[Cat.scala 30:58:@1428.4]
  wire [255:0] _T_1668; // @[Cat.scala 30:58:@1429.4]
  wire [511:0] dat_rsp_pad_value; // @[Cat.scala 30:58:@1430.4]
  wire [511:0] dat_rsp_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1021:23:@1431.4]
  wire [511:0] dat_rsp_l1c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1022:23:@1432.4]
  wire [511:0] dat_rsp_l2c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1023:23:@1433.4]
  wire [511:0] dat_rsp_l3c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1024:23:@1434.4]
  wire [511:0] dat_rsp_l0c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:23:@1435.4]
  wire [511:0] dat_rsp_l1c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1027:23:@1436.4]
  wire [511:0] dat_rsp_l2c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1028:23:@1437.4]
  wire [511:0] dat_rsp_l3c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1029:23:@1438.4]
  wire  _T_1670; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:42:@1440.4]
  wire  _T_1671; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:58:@1441.4]
  wire  _T_1672; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:47:@1442.4]
  wire  _T_1675; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:43:@1443.4]
  wire  _T_1676; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:87:@1444.4]
  wire  _T_1678; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:91:@1445.4]
  wire  _T_1679; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:72:@1446.4]
  wire [255:0] _T_1681; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:171:@1447.4]
  wire [511:0] _T_1682; // @[Cat.scala 30:58:@1448.4]
  wire  _T_1688; // @[NV_NVDLA_CSC_dl_for_check.scala 1041:72:@1452.4]
  wire [255:0] _T_1690; // @[NV_NVDLA_CSC_dl_for_check.scala 1041:171:@1453.4]
  wire [511:0] _T_1691; // @[Cat.scala 30:58:@1454.4]
  wire [511:0] _T_1692; // @[NV_NVDLA_CSC_dl_for_check.scala 1041:27:@1455.4]
  wire [511:0] _T_1693; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:27:@1456.4]
  wire [511:0] dat_rsp_conv_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:27:@1457.4]
  wire [7:0] dat_rsp_conv_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1460.4]
  wire [7:0] dat_rsp_conv_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1462.4]
  wire [7:0] dat_rsp_conv_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1464.4]
  wire [7:0] dat_rsp_conv_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1466.4]
  wire [7:0] dat_rsp_conv_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1468.4]
  wire [7:0] dat_rsp_conv_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1470.4]
  wire [7:0] dat_rsp_conv_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1472.4]
  wire [7:0] dat_rsp_conv_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1474.4]
  wire [7:0] dat_rsp_conv_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1476.4]
  wire [7:0] dat_rsp_conv_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1478.4]
  wire [7:0] dat_rsp_conv_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1480.4]
  wire [7:0] dat_rsp_conv_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1482.4]
  wire [7:0] dat_rsp_conv_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1484.4]
  wire [7:0] dat_rsp_conv_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1486.4]
  wire [7:0] dat_rsp_conv_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1488.4]
  wire [7:0] dat_rsp_conv_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1490.4]
  wire [7:0] dat_rsp_conv_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1492.4]
  wire [7:0] dat_rsp_conv_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1494.4]
  wire [7:0] dat_rsp_conv_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1496.4]
  wire [7:0] dat_rsp_conv_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1498.4]
  wire [7:0] dat_rsp_conv_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1500.4]
  wire [7:0] dat_rsp_conv_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1502.4]
  wire [7:0] dat_rsp_conv_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1504.4]
  wire [7:0] dat_rsp_conv_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1506.4]
  wire [7:0] dat_rsp_conv_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1508.4]
  wire [7:0] dat_rsp_conv_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1510.4]
  wire [7:0] dat_rsp_conv_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1512.4]
  wire [7:0] dat_rsp_conv_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1514.4]
  wire [7:0] dat_rsp_conv_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1516.4]
  wire [7:0] dat_rsp_conv_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1518.4]
  wire [7:0] dat_rsp_conv_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1520.4]
  wire [7:0] dat_rsp_conv_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1522.4]
  wire [7:0] dat_rsp_conv_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1524.4]
  wire [7:0] dat_rsp_conv_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1526.4]
  wire [7:0] dat_rsp_conv_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1528.4]
  wire [7:0] dat_rsp_conv_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1530.4]
  wire [7:0] dat_rsp_conv_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1532.4]
  wire [7:0] dat_rsp_conv_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1534.4]
  wire [7:0] dat_rsp_conv_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1536.4]
  wire [7:0] dat_rsp_conv_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1538.4]
  wire [7:0] dat_rsp_conv_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1540.4]
  wire [7:0] dat_rsp_conv_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1542.4]
  wire [7:0] dat_rsp_conv_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1544.4]
  wire [7:0] dat_rsp_conv_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1546.4]
  wire [7:0] dat_rsp_conv_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1548.4]
  wire [7:0] dat_rsp_conv_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1550.4]
  wire [7:0] dat_rsp_conv_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1552.4]
  wire [7:0] dat_rsp_conv_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1554.4]
  wire [7:0] dat_rsp_conv_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1556.4]
  wire [7:0] dat_rsp_conv_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1558.4]
  wire [7:0] dat_rsp_conv_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1560.4]
  wire [7:0] dat_rsp_conv_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1562.4]
  wire [7:0] dat_rsp_conv_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1564.4]
  wire [7:0] dat_rsp_conv_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1566.4]
  wire [7:0] dat_rsp_conv_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1568.4]
  wire [7:0] dat_rsp_conv_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1570.4]
  wire [7:0] dat_rsp_conv_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1572.4]
  wire [7:0] dat_rsp_conv_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1574.4]
  wire [7:0] dat_rsp_conv_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1576.4]
  wire [7:0] dat_rsp_conv_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1578.4]
  wire [7:0] dat_rsp_conv_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1580.4]
  wire [7:0] dat_rsp_conv_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1582.4]
  wire [7:0] dat_rsp_conv_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1584.4]
  wire [7:0] dat_rsp_conv_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1586.4]
  reg [255:0] dat_rsp_l0_sft_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 1061:28:@1588.4]
  reg [255:0] _RAND_186;
  reg [127:0] dat_rsp_l0_sft_d2; // @[NV_NVDLA_CSC_dl_for_check.scala 1062:28:@1589.4]
  reg [127:0] _RAND_187;
  reg [127:0] dat_rsp_l0_sft_d3; // @[NV_NVDLA_CSC_dl_for_check.scala 1063:28:@1590.4]
  reg [127:0] _RAND_188;
  reg [127:0] dat_rsp_l1_sft_d2; // @[NV_NVDLA_CSC_dl_for_check.scala 1065:28:@1591.4]
  reg [127:0] _RAND_189;
  reg [127:0] dat_rsp_l1_sft_d3; // @[NV_NVDLA_CSC_dl_for_check.scala 1066:28:@1592.4]
  reg [127:0] _RAND_190;
  reg [127:0] dat_rsp_l2_sft_d3; // @[NV_NVDLA_CSC_dl_for_check.scala 1068:28:@1593.4]
  reg [127:0] _RAND_191;
  wire  _T_1834; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:39:@1594.4]
  wire  _T_1835; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:29:@1595.4]
  wire [1023:0] _T_1837; // @[Cat.scala 30:58:@1596.4]
  wire [1023:0] dat_rsp_l0_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:28:@1597.4]
  wire  _T_1838; // @[NV_NVDLA_CSC_dl_for_check.scala 1071:39:@1598.4]
  wire  _T_1839; // @[NV_NVDLA_CSC_dl_for_check.scala 1071:29:@1599.4]
  wire [1023:0] _T_1841; // @[Cat.scala 30:58:@1600.4]
  wire [1023:0] dat_rsp_l1_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1071:28:@1601.4]
  wire  _T_1842; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:39:@1602.4]
  wire  _T_1843; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:29:@1603.4]
  wire [1023:0] _T_1845; // @[Cat.scala 30:58:@1604.4]
  wire [1023:0] dat_rsp_l2_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:28:@1605.4]
  wire  _T_1846; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:39:@1606.4]
  wire  _T_1847; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:29:@1607.4]
  wire [1023:0] _T_1849; // @[Cat.scala 30:58:@1608.4]
  wire [1023:0] dat_rsp_l3_sft_in; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:28:@1609.4]
  wire [10:0] _T_1851; // @[Cat.scala 30:58:@1610.4]
  wire [1023:0] _T_1852; // @[NV_NVDLA_CSC_dl_for_check.scala 1075:41:@1611.4]
  wire [511:0] dat_rsp_l0_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1075:82:@1612.4]
  wire [10:0] _T_1854; // @[Cat.scala 30:58:@1613.4]
  wire [1023:0] _T_1855; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:41:@1614.4]
  wire [511:0] dat_rsp_l1_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:82:@1615.4]
  wire [10:0] _T_1857; // @[Cat.scala 30:58:@1616.4]
  wire [1023:0] _T_1858; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:41:@1617.4]
  wire [511:0] dat_rsp_l2_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:82:@1618.4]
  wire [10:0] _T_1860; // @[Cat.scala 30:58:@1619.4]
  wire [1023:0] _T_1861; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:41:@1620.4]
  wire [511:0] dat_rsp_l3_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:82:@1621.4]
  wire  _T_1862; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:36:@1622.4]
  wire  _T_1863; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:26:@1623.4]
  wire  _T_1866; // @[NV_NVDLA_CSC_dl_for_check.scala 1081:41:@1624.4]
  wire [127:0] _T_1867; // @[NV_NVDLA_CSC_dl_for_check.scala 1081:81:@1625.4]
  wire [511:0] _T_1873; // @[Cat.scala 30:58:@1631.4]
  wire  _T_1875; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:41:@1632.4]
  wire [255:0] _T_1876; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:81:@1633.4]
  wire [511:0] _T_1878; // @[Cat.scala 30:58:@1635.4]
  wire [511:0] _T_1880; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:25:@1637.4]
  wire [511:0] _T_1881; // @[NV_NVDLA_CSC_dl_for_check.scala 1081:25:@1638.4]
  wire [511:0] dat_rsp_img_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:25:@1639.4]
  wire [7:0] dat_rsp_img_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1641.4]
  wire [7:0] dat_rsp_img_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1643.4]
  wire [7:0] dat_rsp_img_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1645.4]
  wire [7:0] dat_rsp_img_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1647.4]
  wire [7:0] dat_rsp_img_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1649.4]
  wire [7:0] dat_rsp_img_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1651.4]
  wire [7:0] dat_rsp_img_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1653.4]
  wire [7:0] dat_rsp_img_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1655.4]
  wire [7:0] dat_rsp_img_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1657.4]
  wire [7:0] dat_rsp_img_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1659.4]
  wire [7:0] dat_rsp_img_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1661.4]
  wire [7:0] dat_rsp_img_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1663.4]
  wire [7:0] dat_rsp_img_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1665.4]
  wire [7:0] dat_rsp_img_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1667.4]
  wire [7:0] dat_rsp_img_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1669.4]
  wire [7:0] dat_rsp_img_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1671.4]
  wire [7:0] dat_rsp_img_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1673.4]
  wire [7:0] dat_rsp_img_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1675.4]
  wire [7:0] dat_rsp_img_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1677.4]
  wire [7:0] dat_rsp_img_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1679.4]
  wire [7:0] dat_rsp_img_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1681.4]
  wire [7:0] dat_rsp_img_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1683.4]
  wire [7:0] dat_rsp_img_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1685.4]
  wire [7:0] dat_rsp_img_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1687.4]
  wire [7:0] dat_rsp_img_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1689.4]
  wire [7:0] dat_rsp_img_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1691.4]
  wire [7:0] dat_rsp_img_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1693.4]
  wire [7:0] dat_rsp_img_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1695.4]
  wire [7:0] dat_rsp_img_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1697.4]
  wire [7:0] dat_rsp_img_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1699.4]
  wire [7:0] dat_rsp_img_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1701.4]
  wire [7:0] dat_rsp_img_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1703.4]
  wire [7:0] dat_rsp_img_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1705.4]
  wire [7:0] dat_rsp_img_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1707.4]
  wire [7:0] dat_rsp_img_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1709.4]
  wire [7:0] dat_rsp_img_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1711.4]
  wire [7:0] dat_rsp_img_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1713.4]
  wire [7:0] dat_rsp_img_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1715.4]
  wire [7:0] dat_rsp_img_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1717.4]
  wire [7:0] dat_rsp_img_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1719.4]
  wire [7:0] dat_rsp_img_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1721.4]
  wire [7:0] dat_rsp_img_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1723.4]
  wire [7:0] dat_rsp_img_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1725.4]
  wire [7:0] dat_rsp_img_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1727.4]
  wire [7:0] dat_rsp_img_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1729.4]
  wire [7:0] dat_rsp_img_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1731.4]
  wire [7:0] dat_rsp_img_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1733.4]
  wire [7:0] dat_rsp_img_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1735.4]
  wire [7:0] dat_rsp_img_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1737.4]
  wire [7:0] dat_rsp_img_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1739.4]
  wire [7:0] dat_rsp_img_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1741.4]
  wire [7:0] dat_rsp_img_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1743.4]
  wire [7:0] dat_rsp_img_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1745.4]
  wire [7:0] dat_rsp_img_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1747.4]
  wire [7:0] dat_rsp_img_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1749.4]
  wire [7:0] dat_rsp_img_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1751.4]
  wire [7:0] dat_rsp_img_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1753.4]
  wire [7:0] dat_rsp_img_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1755.4]
  wire [7:0] dat_rsp_img_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1757.4]
  wire [7:0] dat_rsp_img_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1759.4]
  wire [7:0] dat_rsp_img_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1761.4]
  wire [7:0] dat_rsp_img_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1763.4]
  wire [7:0] dat_rsp_img_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1765.4]
  wire [7:0] dat_rsp_img_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1767.4]
  wire  _T_2016; // @[NV_NVDLA_CSC_dl_for_check.scala 1091:59:@1769.4]
  wire  dat_rsp_sft_d1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1091:41:@1770.4]
  wire  _T_2018; // @[NV_NVDLA_CSC_dl_for_check.scala 1092:59:@1771.4]
  wire  dat_rsp_sft_d2_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1092:41:@1772.4]
  wire  dat_rsp_sft_d3_en; // @[NV_NVDLA_CSC_dl_for_check.scala 1093:41:@1774.4]
  wire [511:0] _GEN_154; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:24:@1775.4]
  wire [255:0] _GEN_155; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:24:@1778.4]
  wire [511:0] _GEN_156; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:24:@1778.4]
  wire [511:0] _GEN_159; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:24:@1782.4]
  wire [318:0] _T_2026; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:55:@1788.4]
  wire [318:0] dat_rsp_ori_mask; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:24:@1789.4]
  wire  _T_2028; // @[NV_NVDLA_CSC_dl_for_check.scala 1113:51:@1790.4]
  wire [63:0] dat_rsp_cur_h_mask_p1; // @[NV_NVDLA_CSC_dl_for_check.scala 1113:32:@1792.4]
  wire  _T_2036; // @[NV_NVDLA_CSC_dl_for_check.scala 1114:51:@1793.4]
  wire [31:0] dat_rsp_cur_h_mask_p2; // @[NV_NVDLA_CSC_dl_for_check.scala 1114:32:@1795.4]
  wire  _T_2044; // @[NV_NVDLA_CSC_dl_for_check.scala 1115:51:@1796.4]
  wire [31:0] dat_rsp_cur_h_mask_p3; // @[NV_NVDLA_CSC_dl_for_check.scala 1115:32:@1798.4]
  wire [31:0] _T_2051; // @[NV_NVDLA_CSC_dl_for_check.scala 1117:57:@1799.4]
  wire [63:0] dat_rsp_cur_h_e2_mask_8b; // @[Cat.scala 30:58:@1801.4]
  wire [15:0] _T_2057; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:57:@1802.4]
  wire [15:0] _T_2058; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:106:@1803.4]
  wire [15:0] _T_2059; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:155:@1804.4]
  wire [63:0] dat_rsp_cur_h_e4_mask_8b; // @[Cat.scala 30:58:@1808.4]
  wire  _T_2068; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:43:@1809.4]
  wire [15:0] _T_2069; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:89:@1810.4]
  wire [63:0] _T_2071; // @[Cat.scala 30:58:@1812.4]
  wire [63:0] _T_2072; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:116:@1813.4]
  wire  _T_2074; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:43:@1814.4]
  wire [31:0] _T_2075; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:89:@1815.4]
  wire [63:0] _T_2076; // @[Cat.scala 30:58:@1816.4]
  wire [63:0] _T_2077; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:116:@1817.4]
  wire [63:0] _T_2078; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:39:@1818.4]
  wire [63:0] _T_2079; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:26:@1819.4]
  wire [63:0] dat_rsp_mask_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:26:@1820.4]
  wire  _T_2080; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:35:@1821.4]
  wire [7:0] dat_rsp_data_w_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire [7:0] dat_rsp_data_w_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  wire  dat_rsp_mask_val_int8_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1823.4]
  wire  dat_rsp_mask_val_int8_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1824.4]
  wire  dat_rsp_mask_val_int8_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1825.4]
  wire  dat_rsp_mask_val_int8_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1826.4]
  wire  dat_rsp_mask_val_int8_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1827.4]
  wire  dat_rsp_mask_val_int8_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1828.4]
  wire  dat_rsp_mask_val_int8_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1829.4]
  wire  dat_rsp_mask_val_int8_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1830.4]
  wire  dat_rsp_mask_val_int8_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1831.4]
  wire  dat_rsp_mask_val_int8_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1832.4]
  wire  dat_rsp_mask_val_int8_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1833.4]
  wire  dat_rsp_mask_val_int8_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1834.4]
  wire  dat_rsp_mask_val_int8_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1835.4]
  wire  dat_rsp_mask_val_int8_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1836.4]
  wire  dat_rsp_mask_val_int8_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1837.4]
  wire  dat_rsp_mask_val_int8_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1838.4]
  wire  dat_rsp_mask_val_int8_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1839.4]
  wire  dat_rsp_mask_val_int8_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1840.4]
  wire  dat_rsp_mask_val_int8_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1841.4]
  wire  dat_rsp_mask_val_int8_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1842.4]
  wire  dat_rsp_mask_val_int8_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1843.4]
  wire  dat_rsp_mask_val_int8_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1844.4]
  wire  dat_rsp_mask_val_int8_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1845.4]
  wire  dat_rsp_mask_val_int8_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1846.4]
  wire  dat_rsp_mask_val_int8_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1847.4]
  wire  dat_rsp_mask_val_int8_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1848.4]
  wire  dat_rsp_mask_val_int8_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1849.4]
  wire  dat_rsp_mask_val_int8_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1850.4]
  wire  dat_rsp_mask_val_int8_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1851.4]
  wire  dat_rsp_mask_val_int8_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1852.4]
  wire  dat_rsp_mask_val_int8_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1853.4]
  wire  dat_rsp_mask_val_int8_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1854.4]
  wire  dat_rsp_mask_val_int8_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1855.4]
  wire  dat_rsp_mask_val_int8_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1856.4]
  wire  dat_rsp_mask_val_int8_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1857.4]
  wire  dat_rsp_mask_val_int8_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1858.4]
  wire  dat_rsp_mask_val_int8_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1859.4]
  wire  dat_rsp_mask_val_int8_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1860.4]
  wire  dat_rsp_mask_val_int8_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1861.4]
  wire  dat_rsp_mask_val_int8_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1862.4]
  wire  dat_rsp_mask_val_int8_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1863.4]
  wire  dat_rsp_mask_val_int8_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1864.4]
  wire  dat_rsp_mask_val_int8_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1865.4]
  wire  dat_rsp_mask_val_int8_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1866.4]
  wire  dat_rsp_mask_val_int8_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1867.4]
  wire  dat_rsp_mask_val_int8_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1868.4]
  wire  dat_rsp_mask_val_int8_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1869.4]
  wire  dat_rsp_mask_val_int8_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1870.4]
  wire  dat_rsp_mask_val_int8_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1871.4]
  wire  dat_rsp_mask_val_int8_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1872.4]
  wire  dat_rsp_mask_val_int8_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1873.4]
  wire  dat_rsp_mask_val_int8_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1874.4]
  wire  dat_rsp_mask_val_int8_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1875.4]
  wire  dat_rsp_mask_val_int8_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1876.4]
  wire  dat_rsp_mask_val_int8_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1877.4]
  wire  dat_rsp_mask_val_int8_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1878.4]
  wire  dat_rsp_mask_val_int8_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1879.4]
  wire  dat_rsp_mask_val_int8_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1880.4]
  wire  dat_rsp_mask_val_int8_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1881.4]
  wire  dat_rsp_mask_val_int8_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1882.4]
  wire  dat_rsp_mask_val_int8_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1883.4]
  wire  dat_rsp_mask_val_int8_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1884.4]
  wire  dat_rsp_mask_val_int8_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1885.4]
  wire  dat_rsp_mask_val_int8_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1886.4]
  wire  _T_2409; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1952.4]
  wire  dat_rsp_mask_w_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1953.4]
  wire  _T_2411; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1954.4]
  wire  dat_rsp_mask_w_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1955.4]
  wire  _T_2413; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1956.4]
  wire  dat_rsp_mask_w_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1957.4]
  wire  _T_2415; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1958.4]
  wire  dat_rsp_mask_w_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1959.4]
  wire  _T_2417; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1960.4]
  wire  dat_rsp_mask_w_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1961.4]
  wire  _T_2419; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1962.4]
  wire  dat_rsp_mask_w_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1963.4]
  wire  _T_2421; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1964.4]
  wire  dat_rsp_mask_w_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1965.4]
  wire  _T_2423; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1966.4]
  wire  dat_rsp_mask_w_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1967.4]
  wire  _T_2425; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1968.4]
  wire  dat_rsp_mask_w_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1969.4]
  wire  _T_2427; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1970.4]
  wire  dat_rsp_mask_w_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1971.4]
  wire  _T_2429; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1972.4]
  wire  dat_rsp_mask_w_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1973.4]
  wire  _T_2431; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1974.4]
  wire  dat_rsp_mask_w_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1975.4]
  wire  _T_2433; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1976.4]
  wire  dat_rsp_mask_w_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1977.4]
  wire  _T_2435; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1978.4]
  wire  dat_rsp_mask_w_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1979.4]
  wire  _T_2437; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1980.4]
  wire  dat_rsp_mask_w_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1981.4]
  wire  _T_2439; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1982.4]
  wire  dat_rsp_mask_w_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1983.4]
  wire  _T_2441; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1984.4]
  wire  dat_rsp_mask_w_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1985.4]
  wire  _T_2443; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1986.4]
  wire  dat_rsp_mask_w_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1987.4]
  wire  _T_2445; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1988.4]
  wire  dat_rsp_mask_w_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1989.4]
  wire  _T_2447; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1990.4]
  wire  dat_rsp_mask_w_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1991.4]
  wire  _T_2449; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1992.4]
  wire  dat_rsp_mask_w_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1993.4]
  wire  _T_2451; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1994.4]
  wire  dat_rsp_mask_w_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1995.4]
  wire  _T_2453; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1996.4]
  wire  dat_rsp_mask_w_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1997.4]
  wire  _T_2455; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1998.4]
  wire  dat_rsp_mask_w_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1999.4]
  wire  _T_2457; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2000.4]
  wire  dat_rsp_mask_w_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2001.4]
  wire  _T_2459; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2002.4]
  wire  dat_rsp_mask_w_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2003.4]
  wire  _T_2461; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2004.4]
  wire  dat_rsp_mask_w_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2005.4]
  wire  _T_2463; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2006.4]
  wire  dat_rsp_mask_w_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2007.4]
  wire  _T_2465; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2008.4]
  wire  dat_rsp_mask_w_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2009.4]
  wire  _T_2467; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2010.4]
  wire  dat_rsp_mask_w_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2011.4]
  wire  _T_2469; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2012.4]
  wire  dat_rsp_mask_w_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2013.4]
  wire  _T_2471; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2014.4]
  wire  dat_rsp_mask_w_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2015.4]
  wire  _T_2473; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2016.4]
  wire  dat_rsp_mask_w_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2017.4]
  wire  _T_2475; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2018.4]
  wire  dat_rsp_mask_w_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2019.4]
  wire  _T_2477; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2020.4]
  wire  dat_rsp_mask_w_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2021.4]
  wire  _T_2479; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2022.4]
  wire  dat_rsp_mask_w_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2023.4]
  wire  _T_2481; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2024.4]
  wire  dat_rsp_mask_w_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2025.4]
  wire  _T_2483; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2026.4]
  wire  dat_rsp_mask_w_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2027.4]
  wire  _T_2485; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2028.4]
  wire  dat_rsp_mask_w_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2029.4]
  wire  _T_2487; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2030.4]
  wire  dat_rsp_mask_w_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2031.4]
  wire  _T_2489; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2032.4]
  wire  dat_rsp_mask_w_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2033.4]
  wire  _T_2491; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2034.4]
  wire  dat_rsp_mask_w_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2035.4]
  wire  _T_2493; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2036.4]
  wire  dat_rsp_mask_w_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2037.4]
  wire  _T_2495; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2038.4]
  wire  dat_rsp_mask_w_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2039.4]
  wire  _T_2497; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2040.4]
  wire  dat_rsp_mask_w_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2041.4]
  wire  _T_2499; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2042.4]
  wire  dat_rsp_mask_w_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2043.4]
  wire  _T_2501; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2044.4]
  wire  dat_rsp_mask_w_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2045.4]
  wire  _T_2503; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2046.4]
  wire  dat_rsp_mask_w_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2047.4]
  wire  _T_2505; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2048.4]
  wire  dat_rsp_mask_w_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2049.4]
  wire  _T_2507; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2050.4]
  wire  dat_rsp_mask_w_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2051.4]
  wire  _T_2509; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2052.4]
  wire  dat_rsp_mask_w_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2053.4]
  wire  _T_2511; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2054.4]
  wire  dat_rsp_mask_w_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2055.4]
  wire  _T_2513; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2056.4]
  wire  dat_rsp_mask_w_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2057.4]
  wire  _T_2515; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2058.4]
  wire  dat_rsp_mask_w_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2059.4]
  wire  _T_2517; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2060.4]
  wire  dat_rsp_mask_w_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2061.4]
  wire  _T_2519; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2062.4]
  wire  dat_rsp_mask_w_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2063.4]
  wire  _T_2521; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2064.4]
  wire  dat_rsp_mask_w_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2065.4]
  wire  _T_2523; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2066.4]
  wire  dat_rsp_mask_w_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2067.4]
  wire  _T_2525; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2068.4]
  wire  dat_rsp_mask_w_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2069.4]
  wire  _T_2527; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2070.4]
  wire  dat_rsp_mask_w_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2071.4]
  wire  _T_2529; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2072.4]
  wire  dat_rsp_mask_w_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2073.4]
  wire  _T_2531; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2074.4]
  wire  dat_rsp_mask_w_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2075.4]
  wire  _T_2533; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2076.4]
  wire  dat_rsp_mask_w_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2077.4]
  wire  _T_2535; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2078.4]
  wire  dat_rsp_mask_w_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2079.4]
  wire  _T_2606; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:54:@2145.4]
  wire  _T_2607; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:39:@2146.4]
  wire  dat_rsp_p0_vld_w; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:37:@2147.4]
  reg  dat_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1133:27:@2148.4]
  reg [31:0] _RAND_192;
  reg [8:0] dat_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1134:27:@2149.4]
  reg [31:0] _RAND_193;
  reg  dat_out_bypass_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_194;
  reg  dat_out_bypass_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_195;
  reg  dat_out_bypass_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_196;
  reg  dat_out_bypass_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_197;
  reg  dat_out_bypass_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_198;
  reg  dat_out_bypass_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_199;
  reg  dat_out_bypass_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_200;
  reg  dat_out_bypass_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_201;
  reg  dat_out_bypass_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_202;
  reg  dat_out_bypass_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_203;
  reg  dat_out_bypass_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_204;
  reg  dat_out_bypass_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_205;
  reg  dat_out_bypass_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_206;
  reg  dat_out_bypass_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_207;
  reg  dat_out_bypass_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_208;
  reg  dat_out_bypass_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_209;
  reg  dat_out_bypass_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_210;
  reg  dat_out_bypass_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_211;
  reg  dat_out_bypass_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_212;
  reg  dat_out_bypass_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_213;
  reg  dat_out_bypass_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_214;
  reg  dat_out_bypass_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_215;
  reg  dat_out_bypass_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_216;
  reg  dat_out_bypass_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_217;
  reg  dat_out_bypass_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_218;
  reg  dat_out_bypass_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_219;
  reg  dat_out_bypass_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_220;
  reg  dat_out_bypass_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_221;
  reg  dat_out_bypass_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_222;
  reg  dat_out_bypass_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_223;
  reg  dat_out_bypass_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_224;
  reg  dat_out_bypass_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_225;
  reg  dat_out_bypass_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_226;
  reg  dat_out_bypass_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_227;
  reg  dat_out_bypass_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_228;
  reg  dat_out_bypass_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_229;
  reg  dat_out_bypass_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_230;
  reg  dat_out_bypass_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_231;
  reg  dat_out_bypass_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_232;
  reg  dat_out_bypass_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_233;
  reg  dat_out_bypass_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_234;
  reg  dat_out_bypass_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_235;
  reg  dat_out_bypass_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_236;
  reg  dat_out_bypass_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_237;
  reg  dat_out_bypass_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_238;
  reg  dat_out_bypass_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_239;
  reg  dat_out_bypass_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_240;
  reg  dat_out_bypass_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_241;
  reg  dat_out_bypass_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_242;
  reg  dat_out_bypass_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_243;
  reg  dat_out_bypass_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_244;
  reg  dat_out_bypass_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_245;
  reg  dat_out_bypass_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_246;
  reg  dat_out_bypass_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_247;
  reg  dat_out_bypass_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_248;
  reg  dat_out_bypass_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_249;
  reg  dat_out_bypass_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_250;
  reg  dat_out_bypass_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_251;
  reg  dat_out_bypass_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_252;
  reg  dat_out_bypass_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_253;
  reg  dat_out_bypass_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_254;
  reg  dat_out_bypass_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_255;
  reg  dat_out_bypass_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_256;
  reg  dat_out_bypass_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1135:34:@2215.4]
  reg [31:0] _RAND_257;
  reg [7:0] dat_out_bypass_data_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_258;
  reg [7:0] dat_out_bypass_data_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_259;
  reg [7:0] dat_out_bypass_data_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_260;
  reg [7:0] dat_out_bypass_data_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_261;
  reg [7:0] dat_out_bypass_data_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_262;
  reg [7:0] dat_out_bypass_data_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_263;
  reg [7:0] dat_out_bypass_data_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_264;
  reg [7:0] dat_out_bypass_data_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_265;
  reg [7:0] dat_out_bypass_data_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_266;
  reg [7:0] dat_out_bypass_data_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_267;
  reg [7:0] dat_out_bypass_data_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_268;
  reg [7:0] dat_out_bypass_data_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_269;
  reg [7:0] dat_out_bypass_data_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_270;
  reg [7:0] dat_out_bypass_data_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_271;
  reg [7:0] dat_out_bypass_data_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_272;
  reg [7:0] dat_out_bypass_data_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_273;
  reg [7:0] dat_out_bypass_data_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_274;
  reg [7:0] dat_out_bypass_data_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_275;
  reg [7:0] dat_out_bypass_data_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_276;
  reg [7:0] dat_out_bypass_data_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_277;
  reg [7:0] dat_out_bypass_data_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_278;
  reg [7:0] dat_out_bypass_data_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_279;
  reg [7:0] dat_out_bypass_data_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_280;
  reg [7:0] dat_out_bypass_data_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_281;
  reg [7:0] dat_out_bypass_data_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_282;
  reg [7:0] dat_out_bypass_data_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_283;
  reg [7:0] dat_out_bypass_data_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_284;
  reg [7:0] dat_out_bypass_data_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_285;
  reg [7:0] dat_out_bypass_data_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_286;
  reg [7:0] dat_out_bypass_data_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_287;
  reg [7:0] dat_out_bypass_data_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_288;
  reg [7:0] dat_out_bypass_data_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_289;
  reg [7:0] dat_out_bypass_data_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_290;
  reg [7:0] dat_out_bypass_data_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_291;
  reg [7:0] dat_out_bypass_data_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_292;
  reg [7:0] dat_out_bypass_data_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_293;
  reg [7:0] dat_out_bypass_data_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_294;
  reg [7:0] dat_out_bypass_data_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_295;
  reg [7:0] dat_out_bypass_data_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_296;
  reg [7:0] dat_out_bypass_data_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_297;
  reg [7:0] dat_out_bypass_data_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_298;
  reg [7:0] dat_out_bypass_data_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_299;
  reg [7:0] dat_out_bypass_data_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_300;
  reg [7:0] dat_out_bypass_data_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_301;
  reg [7:0] dat_out_bypass_data_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_302;
  reg [7:0] dat_out_bypass_data_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_303;
  reg [7:0] dat_out_bypass_data_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_304;
  reg [7:0] dat_out_bypass_data_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_305;
  reg [7:0] dat_out_bypass_data_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_306;
  reg [7:0] dat_out_bypass_data_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_307;
  reg [7:0] dat_out_bypass_data_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_308;
  reg [7:0] dat_out_bypass_data_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_309;
  reg [7:0] dat_out_bypass_data_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_310;
  reg [7:0] dat_out_bypass_data_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_311;
  reg [7:0] dat_out_bypass_data_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_312;
  reg [7:0] dat_out_bypass_data_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_313;
  reg [7:0] dat_out_bypass_data_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_314;
  reg [7:0] dat_out_bypass_data_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_315;
  reg [7:0] dat_out_bypass_data_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_316;
  reg [7:0] dat_out_bypass_data_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_317;
  reg [7:0] dat_out_bypass_data_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_318;
  reg [7:0] dat_out_bypass_data_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_319;
  reg [7:0] dat_out_bypass_data_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_320;
  reg [7:0] dat_out_bypass_data_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1136:30:@2216.4]
  reg [31:0] _RAND_321;
  reg  _T_3147; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:64:@2218.4]
  reg [31:0] _RAND_322;
  reg  _T_3150; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:64:@2219.4]
  reg [31:0] _RAND_323;
  reg  _T_3153; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:64:@2220.4]
  reg [31:0] _RAND_324;
  reg  _T_3156; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:64:@2221.4]
  reg [31:0] _RAND_325;
  reg  _T_3159; // @[NV_NVDLA_CSC_dl_for_check.scala 1139:64:@2222.4]
  reg [31:0] _RAND_326;
  reg [8:0] _T_3164; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:64:@2224.4]
  reg [31:0] _RAND_327;
  reg [8:0] _T_3167; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:64:@2225.4]
  reg [31:0] _RAND_328;
  reg [8:0] _T_3170; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:64:@2226.4]
  reg [31:0] _RAND_329;
  reg [8:0] _T_3173; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:64:@2227.4]
  reg [31:0] _RAND_330;
  reg [8:0] _T_3176; // @[NV_NVDLA_CSC_dl_for_check.scala 1141:64:@2228.4]
  reg [31:0] _RAND_331;
  wire [8:0] _GEN_160; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2232.4]
  wire [8:0] _GEN_161; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2236.4]
  wire [8:0] _GEN_162; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2240.4]
  wire [8:0] _GEN_163; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2244.4]
  wire [8:0] _GEN_164; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2248.4]
  wire  _T_3177; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:40:@2251.4]
  wire  dat_out_pvld_w; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:25:@2252.4]
  wire  _T_3178; // @[NV_NVDLA_CSC_dl_for_check.scala 1154:40:@2253.4]
  wire [8:0] dat_out_flag_w; // @[NV_NVDLA_CSC_dl_for_check.scala 1154:25:@2254.4]
  wire [8:0] _GEN_165; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:21:@2256.4]
  wire  _GEN_166; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_167; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_168; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_169; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_170; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_171; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_172; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_173; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_174; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_175; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_176; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_177; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_178; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_179; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_180; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_181; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_182; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_183; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_184; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_185; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_186; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_187; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_188; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_189; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_190; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_191; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_192; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_193; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_194; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_195; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_196; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_197; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_198; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_199; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_200; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_201; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_202; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_203; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_204; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_205; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_206; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_207; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_208; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_209; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_210; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_211; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_212; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_213; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_214; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_215; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_216; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_217; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_218; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_219; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_220; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_221; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_222; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_223; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_224; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_225; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_226; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_227; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_228; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _GEN_229; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  wire  _T_3179; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2325.4]
  wire  _T_3180; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2329.4]
  wire  _T_3181; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2333.4]
  wire  _T_3182; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2337.4]
  wire  _T_3183; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2341.4]
  wire  _T_3184; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2345.4]
  wire  _T_3185; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2349.4]
  wire  _T_3186; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2353.4]
  wire  _T_3187; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2357.4]
  wire  _T_3188; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2361.4]
  wire  _T_3189; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2365.4]
  wire  _T_3190; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2369.4]
  wire  _T_3191; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2373.4]
  wire  _T_3192; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2377.4]
  wire  _T_3193; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2381.4]
  wire  _T_3194; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2385.4]
  wire  _T_3195; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2389.4]
  wire  _T_3196; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2393.4]
  wire  _T_3197; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2397.4]
  wire  _T_3198; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2401.4]
  wire  _T_3199; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2405.4]
  wire  _T_3200; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2409.4]
  wire  _T_3201; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2413.4]
  wire  _T_3202; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2417.4]
  wire  _T_3203; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2421.4]
  wire  _T_3204; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2425.4]
  wire  _T_3205; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2429.4]
  wire  _T_3206; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2433.4]
  wire  _T_3207; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2437.4]
  wire  _T_3208; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2441.4]
  wire  _T_3209; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2445.4]
  wire  _T_3210; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2449.4]
  wire  _T_3211; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2453.4]
  wire  _T_3212; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2457.4]
  wire  _T_3213; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2461.4]
  wire  _T_3214; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2465.4]
  wire  _T_3215; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2469.4]
  wire  _T_3216; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2473.4]
  wire  _T_3217; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2477.4]
  wire  _T_3218; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2481.4]
  wire  _T_3219; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2485.4]
  wire  _T_3220; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2489.4]
  wire  _T_3221; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2493.4]
  wire  _T_3222; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2497.4]
  wire  _T_3223; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2501.4]
  wire  _T_3224; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2505.4]
  wire  _T_3225; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2509.4]
  wire  _T_3226; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2513.4]
  wire  _T_3227; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2517.4]
  wire  _T_3228; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2521.4]
  wire  _T_3229; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2525.4]
  wire  _T_3230; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2529.4]
  wire  _T_3231; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2533.4]
  wire  _T_3232; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2537.4]
  wire  _T_3233; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2541.4]
  wire  _T_3234; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2545.4]
  wire  _T_3235; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2549.4]
  wire  _T_3236; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2553.4]
  wire  _T_3237; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2557.4]
  wire  _T_3238; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2561.4]
  wire  _T_3239; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2565.4]
  wire  _T_3240; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2569.4]
  wire  _T_3241; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2573.4]
  wire  _T_3242; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2577.4]
  reg  dl_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1182:26:@2711.4]
  reg [31:0] _RAND_332;
  reg  dl_out_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_333;
  reg  dl_out_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_334;
  reg  dl_out_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_335;
  reg  dl_out_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_336;
  reg  dl_out_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_337;
  reg  dl_out_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_338;
  reg  dl_out_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_339;
  reg  dl_out_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_340;
  reg  dl_out_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_341;
  reg  dl_out_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_342;
  reg  dl_out_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_343;
  reg  dl_out_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_344;
  reg  dl_out_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_345;
  reg  dl_out_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_346;
  reg  dl_out_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_347;
  reg  dl_out_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_348;
  reg  dl_out_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_349;
  reg  dl_out_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_350;
  reg  dl_out_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_351;
  reg  dl_out_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_352;
  reg  dl_out_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_353;
  reg  dl_out_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_354;
  reg  dl_out_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_355;
  reg  dl_out_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_356;
  reg  dl_out_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_357;
  reg  dl_out_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_358;
  reg  dl_out_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_359;
  reg  dl_out_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_360;
  reg  dl_out_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_361;
  reg  dl_out_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_362;
  reg  dl_out_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_363;
  reg  dl_out_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_364;
  reg  dl_out_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_365;
  reg  dl_out_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_366;
  reg  dl_out_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_367;
  reg  dl_out_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_368;
  reg  dl_out_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_369;
  reg  dl_out_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_370;
  reg  dl_out_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_371;
  reg  dl_out_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_372;
  reg  dl_out_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_373;
  reg  dl_out_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_374;
  reg  dl_out_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_375;
  reg  dl_out_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_376;
  reg  dl_out_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_377;
  reg  dl_out_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_378;
  reg  dl_out_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_379;
  reg  dl_out_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_380;
  reg  dl_out_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_381;
  reg  dl_out_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_382;
  reg  dl_out_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_383;
  reg  dl_out_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_384;
  reg  dl_out_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_385;
  reg  dl_out_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_386;
  reg  dl_out_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_387;
  reg  dl_out_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_388;
  reg  dl_out_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_389;
  reg  dl_out_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_390;
  reg  dl_out_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_391;
  reg  dl_out_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_392;
  reg  dl_out_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_393;
  reg  dl_out_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_394;
  reg  dl_out_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_395;
  reg  dl_out_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1183:26:@2777.4]
  reg [31:0] _RAND_396;
  reg [8:0] dl_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1184:26:@2778.4]
  reg [31:0] _RAND_397;
  reg [7:0] dl_out_data_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_398;
  reg [7:0] dl_out_data_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_399;
  reg [7:0] dl_out_data_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_400;
  reg [7:0] dl_out_data_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_401;
  reg [7:0] dl_out_data_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_402;
  reg [7:0] dl_out_data_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_403;
  reg [7:0] dl_out_data_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_404;
  reg [7:0] dl_out_data_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_405;
  reg [7:0] dl_out_data_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_406;
  reg [7:0] dl_out_data_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_407;
  reg [7:0] dl_out_data_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_408;
  reg [7:0] dl_out_data_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_409;
  reg [7:0] dl_out_data_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_410;
  reg [7:0] dl_out_data_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_411;
  reg [7:0] dl_out_data_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_412;
  reg [7:0] dl_out_data_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_413;
  reg [7:0] dl_out_data_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_414;
  reg [7:0] dl_out_data_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_415;
  reg [7:0] dl_out_data_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_416;
  reg [7:0] dl_out_data_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_417;
  reg [7:0] dl_out_data_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_418;
  reg [7:0] dl_out_data_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_419;
  reg [7:0] dl_out_data_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_420;
  reg [7:0] dl_out_data_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_421;
  reg [7:0] dl_out_data_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_422;
  reg [7:0] dl_out_data_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_423;
  reg [7:0] dl_out_data_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_424;
  reg [7:0] dl_out_data_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_425;
  reg [7:0] dl_out_data_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_426;
  reg [7:0] dl_out_data_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_427;
  reg [7:0] dl_out_data_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_428;
  reg [7:0] dl_out_data_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_429;
  reg [7:0] dl_out_data_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_430;
  reg [7:0] dl_out_data_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_431;
  reg [7:0] dl_out_data_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_432;
  reg [7:0] dl_out_data_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_433;
  reg [7:0] dl_out_data_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_434;
  reg [7:0] dl_out_data_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_435;
  reg [7:0] dl_out_data_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_436;
  reg [7:0] dl_out_data_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_437;
  reg [7:0] dl_out_data_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_438;
  reg [7:0] dl_out_data_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_439;
  reg [7:0] dl_out_data_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_440;
  reg [7:0] dl_out_data_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_441;
  reg [7:0] dl_out_data_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_442;
  reg [7:0] dl_out_data_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_443;
  reg [7:0] dl_out_data_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_444;
  reg [7:0] dl_out_data_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_445;
  reg [7:0] dl_out_data_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_446;
  reg [7:0] dl_out_data_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_447;
  reg [7:0] dl_out_data_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_448;
  reg [7:0] dl_out_data_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_449;
  reg [7:0] dl_out_data_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_450;
  reg [7:0] dl_out_data_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_451;
  reg [7:0] dl_out_data_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_452;
  reg [7:0] dl_out_data_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_453;
  reg [7:0] dl_out_data_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_454;
  reg [7:0] dl_out_data_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_455;
  reg [7:0] dl_out_data_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_456;
  reg [7:0] dl_out_data_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_457;
  reg [7:0] dl_out_data_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_458;
  reg [7:0] dl_out_data_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_459;
  reg [7:0] dl_out_data_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_460;
  reg [7:0] dl_out_data_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1185:22:@2779.4]
  reg [31:0] _RAND_461;
  wire  _T_4044; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:38:@2780.4]
  wire [7:0] dat_out_data_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire [7:0] dat_out_data_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  wire  _T_4176; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:24:@2782.4]
  wire  _T_4311; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:38:@2848.4]
  wire  _T_4312_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  _T_4312_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  wire  dat_out_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  dat_out_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  wire  _T_4575; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:19:@2852.4]
  wire  _GEN_294; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_295; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_296; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_297; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_298; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_299; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_300; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_301; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_302; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_303; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_304; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_305; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_306; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_307; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_308; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_309; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_310; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_311; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_312; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_313; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_314; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_315; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_316; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_317; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_318; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_319; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_320; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_321; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_322; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_323; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_324; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_325; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_326; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_327; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_328; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_329; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_330; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_331; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_332; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_333; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_334; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_335; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_336; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_337; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_338; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_339; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_340; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_341; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_342; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_343; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_344; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_345; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_346; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_347; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_348; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_349; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_350; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_351; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_352; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_353; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_354; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_355; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_356; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire  _GEN_357; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  wire [8:0] _GEN_358; // @[NV_NVDLA_CSC_dl_for_check.scala 1195:19:@2919.4]
  reg  dl_out_pvld_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 1208:29:@3114.4]
  reg [31:0] _RAND_462;
  wire  _T_4578; // @[NV_NVDLA_CSC_dl_for_check.scala 1209:27:@3116.4]
  wire [8:0] sc2mac_dat_pd_w; // @[NV_NVDLA_CSC_dl_for_check.scala 1209:26:@3117.4]
  reg  _T_4582; // @[NV_NVDLA_CSC_dl_for_check.scala 1211:32:@3118.4]
  reg [31:0] _RAND_463;
  reg  _T_4585; // @[NV_NVDLA_CSC_dl_for_check.scala 1212:32:@3121.4]
  reg [31:0] _RAND_464;
  wire  _T_4587; // @[NV_NVDLA_CSC_dl_for_check.scala 1213:80:@3124.4]
  reg [8:0] _T_4589; // @[Reg.scala 19:20:@3125.4]
  reg [31:0] _RAND_465;
  wire [8:0] _GEN_423; // @[Reg.scala 20:19:@3126.4]
  reg [8:0] _T_4593; // @[Reg.scala 19:20:@3131.4]
  reg [31:0] _RAND_466;
  wire [8:0] _GEN_424; // @[Reg.scala 20:19:@3132.4]
  reg  _T_4861_0; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_467;
  reg  _T_4861_1; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_468;
  reg  _T_4861_2; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_469;
  reg  _T_4861_3; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_470;
  reg  _T_4861_4; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_471;
  reg  _T_4861_5; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_472;
  reg  _T_4861_6; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_473;
  reg  _T_4861_7; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_474;
  reg  _T_4861_8; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_475;
  reg  _T_4861_9; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_476;
  reg  _T_4861_10; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_477;
  reg  _T_4861_11; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_478;
  reg  _T_4861_12; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_479;
  reg  _T_4861_13; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_480;
  reg  _T_4861_14; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_481;
  reg  _T_4861_15; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_482;
  reg  _T_4861_16; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_483;
  reg  _T_4861_17; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_484;
  reg  _T_4861_18; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_485;
  reg  _T_4861_19; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_486;
  reg  _T_4861_20; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_487;
  reg  _T_4861_21; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_488;
  reg  _T_4861_22; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_489;
  reg  _T_4861_23; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_490;
  reg  _T_4861_24; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_491;
  reg  _T_4861_25; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_492;
  reg  _T_4861_26; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_493;
  reg  _T_4861_27; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_494;
  reg  _T_4861_28; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_495;
  reg  _T_4861_29; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_496;
  reg  _T_4861_30; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_497;
  reg  _T_4861_31; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_498;
  reg  _T_4861_32; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_499;
  reg  _T_4861_33; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_500;
  reg  _T_4861_34; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_501;
  reg  _T_4861_35; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_502;
  reg  _T_4861_36; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_503;
  reg  _T_4861_37; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_504;
  reg  _T_4861_38; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_505;
  reg  _T_4861_39; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_506;
  reg  _T_4861_40; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_507;
  reg  _T_4861_41; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_508;
  reg  _T_4861_42; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_509;
  reg  _T_4861_43; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_510;
  reg  _T_4861_44; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_511;
  reg  _T_4861_45; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_512;
  reg  _T_4861_46; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_513;
  reg  _T_4861_47; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_514;
  reg  _T_4861_48; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_515;
  reg  _T_4861_49; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_516;
  reg  _T_4861_50; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_517;
  reg  _T_4861_51; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_518;
  reg  _T_4861_52; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_519;
  reg  _T_4861_53; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_520;
  reg  _T_4861_54; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_521;
  reg  _T_4861_55; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_522;
  reg  _T_4861_56; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_523;
  reg  _T_4861_57; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_524;
  reg  _T_4861_58; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_525;
  reg  _T_4861_59; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_526;
  reg  _T_4861_60; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_527;
  reg  _T_4861_61; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_528;
  reg  _T_4861_62; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_529;
  reg  _T_4861_63; // @[Reg.scala 19:20:@3202.4]
  reg [31:0] _RAND_530;
  wire  _GEN_425; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_426; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_427; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_428; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_429; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_430; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_431; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_432; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_433; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_434; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_435; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_436; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_437; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_438; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_439; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_440; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_441; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_442; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_443; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_444; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_445; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_446; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_447; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_448; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_449; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_450; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_451; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_452; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_453; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_454; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_455; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_456; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_457; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_458; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_459; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_460; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_461; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_462; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_463; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_464; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_465; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_466; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_467; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_468; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_469; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_470; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_471; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_472; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_473; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_474; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_475; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_476; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_477; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_478; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_479; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_480; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_481; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_482; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_483; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_484; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_485; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_486; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_487; // @[Reg.scala 20:19:@3203.4]
  wire  _GEN_488; // @[Reg.scala 20:19:@3203.4]
  wire [7:0] _T_5064; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3275.4]
  wire [15:0] _T_5072; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3283.4]
  wire [7:0] _T_5079; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3290.4]
  wire [31:0] _T_5088; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3299.4]
  wire [7:0] _T_5095; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3306.4]
  wire [15:0] _T_5103; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3314.4]
  wire [7:0] _T_5110; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3321.4]
  wire [31:0] _T_5119; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3330.4]
  reg  _T_5388_0; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_531;
  reg  _T_5388_1; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_532;
  reg  _T_5388_2; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_533;
  reg  _T_5388_3; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_534;
  reg  _T_5388_4; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_535;
  reg  _T_5388_5; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_536;
  reg  _T_5388_6; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_537;
  reg  _T_5388_7; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_538;
  reg  _T_5388_8; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_539;
  reg  _T_5388_9; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_540;
  reg  _T_5388_10; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_541;
  reg  _T_5388_11; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_542;
  reg  _T_5388_12; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_543;
  reg  _T_5388_13; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_544;
  reg  _T_5388_14; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_545;
  reg  _T_5388_15; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_546;
  reg  _T_5388_16; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_547;
  reg  _T_5388_17; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_548;
  reg  _T_5388_18; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_549;
  reg  _T_5388_19; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_550;
  reg  _T_5388_20; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_551;
  reg  _T_5388_21; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_552;
  reg  _T_5388_22; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_553;
  reg  _T_5388_23; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_554;
  reg  _T_5388_24; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_555;
  reg  _T_5388_25; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_556;
  reg  _T_5388_26; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_557;
  reg  _T_5388_27; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_558;
  reg  _T_5388_28; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_559;
  reg  _T_5388_29; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_560;
  reg  _T_5388_30; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_561;
  reg  _T_5388_31; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_562;
  reg  _T_5388_32; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_563;
  reg  _T_5388_33; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_564;
  reg  _T_5388_34; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_565;
  reg  _T_5388_35; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_566;
  reg  _T_5388_36; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_567;
  reg  _T_5388_37; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_568;
  reg  _T_5388_38; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_569;
  reg  _T_5388_39; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_570;
  reg  _T_5388_40; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_571;
  reg  _T_5388_41; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_572;
  reg  _T_5388_42; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_573;
  reg  _T_5388_43; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_574;
  reg  _T_5388_44; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_575;
  reg  _T_5388_45; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_576;
  reg  _T_5388_46; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_577;
  reg  _T_5388_47; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_578;
  reg  _T_5388_48; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_579;
  reg  _T_5388_49; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_580;
  reg  _T_5388_50; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_581;
  reg  _T_5388_51; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_582;
  reg  _T_5388_52; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_583;
  reg  _T_5388_53; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_584;
  reg  _T_5388_54; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_585;
  reg  _T_5388_55; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_586;
  reg  _T_5388_56; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_587;
  reg  _T_5388_57; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_588;
  reg  _T_5388_58; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_589;
  reg  _T_5388_59; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_590;
  reg  _T_5388_60; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_591;
  reg  _T_5388_61; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_592;
  reg  _T_5388_62; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_593;
  reg  _T_5388_63; // @[Reg.scala 19:20:@3399.4]
  reg [31:0] _RAND_594;
  wire  _GEN_489; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_490; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_491; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_492; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_493; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_494; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_495; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_496; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_497; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_498; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_499; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_500; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_501; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_502; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_503; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_504; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_505; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_506; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_507; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_508; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_509; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_510; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_511; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_512; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_513; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_514; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_515; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_516; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_517; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_518; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_519; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_520; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_521; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_522; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_523; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_524; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_525; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_526; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_527; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_528; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_529; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_530; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_531; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_532; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_533; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_534; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_535; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_536; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_537; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_538; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_539; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_540; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_541; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_542; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_543; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_544; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_545; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_546; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_547; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_548; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_549; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_550; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_551; // @[Reg.scala 20:19:@3400.4]
  wire  _GEN_552; // @[Reg.scala 20:19:@3400.4]
  wire [7:0] _T_5591; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3472.4]
  wire [15:0] _T_5599; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3480.4]
  wire [7:0] _T_5606; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3487.4]
  wire [31:0] _T_5615; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3496.4]
  wire [7:0] _T_5622; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3503.4]
  wire [15:0] _T_5630; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3511.4]
  wire [7:0] _T_5637; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3518.4]
  wire [31:0] _T_5646; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3527.4]
  reg [7:0] _T_5649; // @[Reg.scala 11:16:@3530.4]
  reg [31:0] _RAND_595;
  reg [7:0] _T_5651; // @[Reg.scala 11:16:@3535.4]
  reg [31:0] _RAND_596;
  reg [7:0] _T_5653; // @[Reg.scala 11:16:@3540.4]
  reg [31:0] _RAND_597;
  reg [7:0] _T_5655; // @[Reg.scala 11:16:@3545.4]
  reg [31:0] _RAND_598;
  reg [7:0] _T_5657; // @[Reg.scala 11:16:@3550.4]
  reg [31:0] _RAND_599;
  reg [7:0] _T_5659; // @[Reg.scala 11:16:@3555.4]
  reg [31:0] _RAND_600;
  reg [7:0] _T_5661; // @[Reg.scala 11:16:@3560.4]
  reg [31:0] _RAND_601;
  reg [7:0] _T_5663; // @[Reg.scala 11:16:@3565.4]
  reg [31:0] _RAND_602;
  reg [7:0] _T_5665; // @[Reg.scala 11:16:@3570.4]
  reg [31:0] _RAND_603;
  reg [7:0] _T_5667; // @[Reg.scala 11:16:@3575.4]
  reg [31:0] _RAND_604;
  reg [7:0] _T_5669; // @[Reg.scala 11:16:@3580.4]
  reg [31:0] _RAND_605;
  reg [7:0] _T_5671; // @[Reg.scala 11:16:@3585.4]
  reg [31:0] _RAND_606;
  reg [7:0] _T_5673; // @[Reg.scala 11:16:@3590.4]
  reg [31:0] _RAND_607;
  reg [7:0] _T_5675; // @[Reg.scala 11:16:@3595.4]
  reg [31:0] _RAND_608;
  reg [7:0] _T_5677; // @[Reg.scala 11:16:@3600.4]
  reg [31:0] _RAND_609;
  reg [7:0] _T_5679; // @[Reg.scala 11:16:@3605.4]
  reg [31:0] _RAND_610;
  reg [7:0] _T_5681; // @[Reg.scala 11:16:@3610.4]
  reg [31:0] _RAND_611;
  reg [7:0] _T_5683; // @[Reg.scala 11:16:@3615.4]
  reg [31:0] _RAND_612;
  reg [7:0] _T_5685; // @[Reg.scala 11:16:@3620.4]
  reg [31:0] _RAND_613;
  reg [7:0] _T_5687; // @[Reg.scala 11:16:@3625.4]
  reg [31:0] _RAND_614;
  reg [7:0] _T_5689; // @[Reg.scala 11:16:@3630.4]
  reg [31:0] _RAND_615;
  reg [7:0] _T_5691; // @[Reg.scala 11:16:@3635.4]
  reg [31:0] _RAND_616;
  reg [7:0] _T_5693; // @[Reg.scala 11:16:@3640.4]
  reg [31:0] _RAND_617;
  reg [7:0] _T_5695; // @[Reg.scala 11:16:@3645.4]
  reg [31:0] _RAND_618;
  reg [7:0] _T_5697; // @[Reg.scala 11:16:@3650.4]
  reg [31:0] _RAND_619;
  reg [7:0] _T_5699; // @[Reg.scala 11:16:@3655.4]
  reg [31:0] _RAND_620;
  reg [7:0] _T_5701; // @[Reg.scala 11:16:@3660.4]
  reg [31:0] _RAND_621;
  reg [7:0] _T_5703; // @[Reg.scala 11:16:@3665.4]
  reg [31:0] _RAND_622;
  reg [7:0] _T_5705; // @[Reg.scala 11:16:@3670.4]
  reg [31:0] _RAND_623;
  reg [7:0] _T_5707; // @[Reg.scala 11:16:@3675.4]
  reg [31:0] _RAND_624;
  reg [7:0] _T_5709; // @[Reg.scala 11:16:@3680.4]
  reg [31:0] _RAND_625;
  reg [7:0] _T_5711; // @[Reg.scala 11:16:@3685.4]
  reg [31:0] _RAND_626;
  reg [7:0] _T_5713; // @[Reg.scala 11:16:@3690.4]
  reg [31:0] _RAND_627;
  reg [7:0] _T_5715; // @[Reg.scala 11:16:@3695.4]
  reg [31:0] _RAND_628;
  reg [7:0] _T_5717; // @[Reg.scala 11:16:@3700.4]
  reg [31:0] _RAND_629;
  reg [7:0] _T_5719; // @[Reg.scala 11:16:@3705.4]
  reg [31:0] _RAND_630;
  reg [7:0] _T_5721; // @[Reg.scala 11:16:@3710.4]
  reg [31:0] _RAND_631;
  reg [7:0] _T_5723; // @[Reg.scala 11:16:@3715.4]
  reg [31:0] _RAND_632;
  reg [7:0] _T_5725; // @[Reg.scala 11:16:@3720.4]
  reg [31:0] _RAND_633;
  reg [7:0] _T_5727; // @[Reg.scala 11:16:@3725.4]
  reg [31:0] _RAND_634;
  reg [7:0] _T_5729; // @[Reg.scala 11:16:@3730.4]
  reg [31:0] _RAND_635;
  reg [7:0] _T_5731; // @[Reg.scala 11:16:@3735.4]
  reg [31:0] _RAND_636;
  reg [7:0] _T_5733; // @[Reg.scala 11:16:@3740.4]
  reg [31:0] _RAND_637;
  reg [7:0] _T_5735; // @[Reg.scala 11:16:@3745.4]
  reg [31:0] _RAND_638;
  reg [7:0] _T_5737; // @[Reg.scala 11:16:@3750.4]
  reg [31:0] _RAND_639;
  reg [7:0] _T_5739; // @[Reg.scala 11:16:@3755.4]
  reg [31:0] _RAND_640;
  reg [7:0] _T_5741; // @[Reg.scala 11:16:@3760.4]
  reg [31:0] _RAND_641;
  reg [7:0] _T_5743; // @[Reg.scala 11:16:@3765.4]
  reg [31:0] _RAND_642;
  reg [7:0] _T_5745; // @[Reg.scala 11:16:@3770.4]
  reg [31:0] _RAND_643;
  reg [7:0] _T_5747; // @[Reg.scala 11:16:@3775.4]
  reg [31:0] _RAND_644;
  reg [7:0] _T_5749; // @[Reg.scala 11:16:@3780.4]
  reg [31:0] _RAND_645;
  reg [7:0] _T_5751; // @[Reg.scala 11:16:@3785.4]
  reg [31:0] _RAND_646;
  reg [7:0] _T_5753; // @[Reg.scala 11:16:@3790.4]
  reg [31:0] _RAND_647;
  reg [7:0] _T_5755; // @[Reg.scala 11:16:@3795.4]
  reg [31:0] _RAND_648;
  reg [7:0] _T_5757; // @[Reg.scala 11:16:@3800.4]
  reg [31:0] _RAND_649;
  reg [7:0] _T_5759; // @[Reg.scala 11:16:@3805.4]
  reg [31:0] _RAND_650;
  reg [7:0] _T_5761; // @[Reg.scala 11:16:@3810.4]
  reg [31:0] _RAND_651;
  reg [7:0] _T_5763; // @[Reg.scala 11:16:@3815.4]
  reg [31:0] _RAND_652;
  reg [7:0] _T_5765; // @[Reg.scala 11:16:@3820.4]
  reg [31:0] _RAND_653;
  reg [7:0] _T_5767; // @[Reg.scala 11:16:@3825.4]
  reg [31:0] _RAND_654;
  reg [7:0] _T_5769; // @[Reg.scala 11:16:@3830.4]
  reg [31:0] _RAND_655;
  reg [7:0] _T_5771; // @[Reg.scala 11:16:@3835.4]
  reg [31:0] _RAND_656;
  reg [7:0] _T_5773; // @[Reg.scala 11:16:@3840.4]
  reg [31:0] _RAND_657;
  reg [7:0] _T_5775; // @[Reg.scala 11:16:@3845.4]
  reg [31:0] _RAND_658;
  reg [7:0] _T_5777; // @[Reg.scala 11:16:@3850.4]
  reg [31:0] _RAND_659;
  reg [7:0] _T_5779; // @[Reg.scala 11:16:@3855.4]
  reg [31:0] _RAND_660;
  reg [7:0] _T_5781; // @[Reg.scala 11:16:@3860.4]
  reg [31:0] _RAND_661;
  reg [7:0] _T_5783; // @[Reg.scala 11:16:@3865.4]
  reg [31:0] _RAND_662;
  reg [7:0] _T_5785; // @[Reg.scala 11:16:@3870.4]
  reg [31:0] _RAND_663;
  reg [7:0] _T_5787; // @[Reg.scala 11:16:@3875.4]
  reg [31:0] _RAND_664;
  reg [7:0] _T_5789; // @[Reg.scala 11:16:@3880.4]
  reg [31:0] _RAND_665;
  reg [7:0] _T_5791; // @[Reg.scala 11:16:@3885.4]
  reg [31:0] _RAND_666;
  reg [7:0] _T_5793; // @[Reg.scala 11:16:@3890.4]
  reg [31:0] _RAND_667;
  reg [7:0] _T_5795; // @[Reg.scala 11:16:@3895.4]
  reg [31:0] _RAND_668;
  reg [7:0] _T_5797; // @[Reg.scala 11:16:@3900.4]
  reg [31:0] _RAND_669;
  reg [7:0] _T_5799; // @[Reg.scala 11:16:@3905.4]
  reg [31:0] _RAND_670;
  reg [7:0] _T_5801; // @[Reg.scala 11:16:@3910.4]
  reg [31:0] _RAND_671;
  reg [7:0] _T_5803; // @[Reg.scala 11:16:@3915.4]
  reg [31:0] _RAND_672;
  reg [7:0] _T_5805; // @[Reg.scala 11:16:@3920.4]
  reg [31:0] _RAND_673;
  reg [7:0] _T_5807; // @[Reg.scala 11:16:@3925.4]
  reg [31:0] _RAND_674;
  reg [7:0] _T_5809; // @[Reg.scala 11:16:@3930.4]
  reg [31:0] _RAND_675;
  reg [7:0] _T_5811; // @[Reg.scala 11:16:@3935.4]
  reg [31:0] _RAND_676;
  reg [7:0] _T_5813; // @[Reg.scala 11:16:@3940.4]
  reg [31:0] _RAND_677;
  reg [7:0] _T_5815; // @[Reg.scala 11:16:@3945.4]
  reg [31:0] _RAND_678;
  reg [7:0] _T_5817; // @[Reg.scala 11:16:@3950.4]
  reg [31:0] _RAND_679;
  reg [7:0] _T_5819; // @[Reg.scala 11:16:@3955.4]
  reg [31:0] _RAND_680;
  reg [7:0] _T_5821; // @[Reg.scala 11:16:@3960.4]
  reg [31:0] _RAND_681;
  reg [7:0] _T_5823; // @[Reg.scala 11:16:@3965.4]
  reg [31:0] _RAND_682;
  reg [7:0] _T_5825; // @[Reg.scala 11:16:@3970.4]
  reg [31:0] _RAND_683;
  reg [7:0] _T_5827; // @[Reg.scala 11:16:@3975.4]
  reg [31:0] _RAND_684;
  reg [7:0] _T_5829; // @[Reg.scala 11:16:@3980.4]
  reg [31:0] _RAND_685;
  reg [7:0] _T_5831; // @[Reg.scala 11:16:@3985.4]
  reg [31:0] _RAND_686;
  reg [7:0] _T_5833; // @[Reg.scala 11:16:@3990.4]
  reg [31:0] _RAND_687;
  reg [7:0] _T_5835; // @[Reg.scala 11:16:@3995.4]
  reg [31:0] _RAND_688;
  reg [7:0] _T_5837; // @[Reg.scala 11:16:@4000.4]
  reg [31:0] _RAND_689;
  reg [7:0] _T_5839; // @[Reg.scala 11:16:@4005.4]
  reg [31:0] _RAND_690;
  reg [7:0] _T_5841; // @[Reg.scala 11:16:@4010.4]
  reg [31:0] _RAND_691;
  reg [7:0] _T_5843; // @[Reg.scala 11:16:@4015.4]
  reg [31:0] _RAND_692;
  reg [7:0] _T_5845; // @[Reg.scala 11:16:@4020.4]
  reg [31:0] _RAND_693;
  reg [7:0] _T_5847; // @[Reg.scala 11:16:@4025.4]
  reg [31:0] _RAND_694;
  reg [7:0] _T_5849; // @[Reg.scala 11:16:@4030.4]
  reg [31:0] _RAND_695;
  reg [7:0] _T_5851; // @[Reg.scala 11:16:@4035.4]
  reg [31:0] _RAND_696;
  reg [7:0] _T_5853; // @[Reg.scala 11:16:@4040.4]
  reg [31:0] _RAND_697;
  reg [7:0] _T_5855; // @[Reg.scala 11:16:@4045.4]
  reg [31:0] _RAND_698;
  reg [7:0] _T_5857; // @[Reg.scala 11:16:@4050.4]
  reg [31:0] _RAND_699;
  reg [7:0] _T_5859; // @[Reg.scala 11:16:@4055.4]
  reg [31:0] _RAND_700;
  reg [7:0] _T_5861; // @[Reg.scala 11:16:@4060.4]
  reg [31:0] _RAND_701;
  reg [7:0] _T_5863; // @[Reg.scala 11:16:@4065.4]
  reg [31:0] _RAND_702;
  reg [7:0] _T_5865; // @[Reg.scala 11:16:@4070.4]
  reg [31:0] _RAND_703;
  reg [7:0] _T_5867; // @[Reg.scala 11:16:@4075.4]
  reg [31:0] _RAND_704;
  reg [7:0] _T_5869; // @[Reg.scala 11:16:@4080.4]
  reg [31:0] _RAND_705;
  reg [7:0] _T_5871; // @[Reg.scala 11:16:@4085.4]
  reg [31:0] _RAND_706;
  reg [7:0] _T_5873; // @[Reg.scala 11:16:@4090.4]
  reg [31:0] _RAND_707;
  reg [7:0] _T_5875; // @[Reg.scala 11:16:@4095.4]
  reg [31:0] _RAND_708;
  reg [7:0] _T_5877; // @[Reg.scala 11:16:@4100.4]
  reg [31:0] _RAND_709;
  reg [7:0] _T_5879; // @[Reg.scala 11:16:@4105.4]
  reg [31:0] _RAND_710;
  reg [7:0] _T_5881; // @[Reg.scala 11:16:@4110.4]
  reg [31:0] _RAND_711;
  reg [7:0] _T_5883; // @[Reg.scala 11:16:@4115.4]
  reg [31:0] _RAND_712;
  reg [7:0] _T_5885; // @[Reg.scala 11:16:@4120.4]
  reg [31:0] _RAND_713;
  reg [7:0] _T_5887; // @[Reg.scala 11:16:@4125.4]
  reg [31:0] _RAND_714;
  reg [7:0] _T_5889; // @[Reg.scala 11:16:@4130.4]
  reg [31:0] _RAND_715;
  reg [7:0] _T_5891; // @[Reg.scala 11:16:@4135.4]
  reg [31:0] _RAND_716;
  reg [7:0] _T_5893; // @[Reg.scala 11:16:@4140.4]
  reg [31:0] _RAND_717;
  reg [7:0] _T_5895; // @[Reg.scala 11:16:@4145.4]
  reg [31:0] _RAND_718;
  reg [7:0] _T_5897; // @[Reg.scala 11:16:@4150.4]
  reg [31:0] _RAND_719;
  reg [7:0] _T_5899; // @[Reg.scala 11:16:@4155.4]
  reg [31:0] _RAND_720;
  reg [7:0] _T_5901; // @[Reg.scala 11:16:@4160.4]
  reg [31:0] _RAND_721;
  reg [7:0] _T_5903; // @[Reg.scala 11:16:@4165.4]
  reg [31:0] _RAND_722;
  assign _T_207 = io_nvdla_core_rstn == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 81:38:@8.4]
  assign is_sg_idle = io_sc_state == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 85:31:@9.4]
  assign is_sg_done = io_sc_state == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 87:31:@11.4]
  assign layer_st = io_reg2dp_op_en & is_sg_idle; // @[NV_NVDLA_CSC_dl_for_check.scala 94:32:@14.4]
  assign is_conv = io_reg2dp_conv_mode == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 96:35:@16.4]
  assign is_img = is_conv & io_reg2dp_datain_format; // @[NV_NVDLA_CSC_dl_for_check.scala 97:22:@17.4]
  assign _T_216 = 7'h9 << io_reg2dp_y_extension; // @[NV_NVDLA_CSC_dl_for_check.scala 105:53:@18.4]
  assign _T_218 = is_img ? _T_216 : 7'h8; // @[NV_NVDLA_CSC_dl_for_check.scala 105:24:@19.4]
  assign sub_h_total_w = _T_218[5:3]; // @[NV_NVDLA_CSC_dl_for_check.scala 105:100:@20.4]
  assign sub_h_cmp_w = is_img ? sub_h_total_w : 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 106:22:@21.4]
  assign _T_221 = sub_h_cmp_w - 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 107:34:@22.4]
  assign dataout_w_init = $unsigned(_T_221); // @[NV_NVDLA_CSC_dl_for_check.scala 107:34:@23.4]
  assign conv_x_stride_w = io_reg2dp_conv_x_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 108:73:@24.4]
  assign _T_225 = io_reg2dp_datain_channel_ext[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 109:62:@26.4]
  assign _T_228 = {conv_x_stride_w,2'h0}; // @[Cat.scala 30:58:@27.4]
  assign _T_231 = {conv_x_stride_w,1'h0}; // @[Cat.scala 30:58:@28.4]
  assign _GEN_681 = {{1'd0}, conv_x_stride_w}; // @[NV_NVDLA_CSC_dl_for_check.scala 111:74:@29.4]
  assign _T_232 = _T_231 + _GEN_681; // @[NV_NVDLA_CSC_dl_for_check.scala 111:74:@29.4]
  assign _T_233 = 2'h2 == _T_225; // @[Mux.scala 46:19:@30.4]
  assign _T_234 = _T_233 ? _T_232 : {{2'd0}, conv_x_stride_w}; // @[Mux.scala 46:16:@31.4]
  assign _T_235 = 2'h3 == _T_225; // @[Mux.scala 46:19:@32.4]
  assign pixel_x_stride_w = _T_235 ? _T_228 : _T_234; // @[Mux.scala 46:16:@33.4]
  assign _T_237 = io_reg2dp_weight_channel_ext >= 13'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 113:88:@34.4]
  assign _T_243 = io_reg2dp_weight_channel_ext[5:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 113:172:@36.4]
  assign _T_244 = _T_237 ? 6'h3f : _T_243; // @[NV_NVDLA_CSC_dl_for_check.scala 113:58:@37.4]
  assign _T_247 = {pixel_x_stride_w,1'h0}; // @[Cat.scala 30:58:@38.4]
  assign _GEN_682 = {{1'd0}, pixel_x_stride_w}; // @[NV_NVDLA_CSC_dl_for_check.scala 114:81:@39.4]
  assign _T_248 = _T_247 + _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 114:81:@39.4]
  assign _T_249 = _T_247 + _GEN_682; // @[NV_NVDLA_CSC_dl_for_check.scala 114:81:@40.4]
  assign _GEN_683 = {{1'd0}, _T_243}; // @[NV_NVDLA_CSC_dl_for_check.scala 114:100:@42.4]
  assign _T_251 = _T_249 + _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 114:100:@42.4]
  assign _T_252 = _T_249 + _GEN_683; // @[NV_NVDLA_CSC_dl_for_check.scala 114:100:@43.4]
  assign _T_255 = pixel_x_stride_w + _T_243; // @[NV_NVDLA_CSC_dl_for_check.scala 115:58:@45.4]
  assign _T_256 = pixel_x_stride_w + _T_243; // @[NV_NVDLA_CSC_dl_for_check.scala 115:58:@46.4]
  assign _T_257 = 2'h1 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@47.4]
  assign _T_258 = _T_257 ? _T_256 : _T_244; // @[Mux.scala 46:16:@48.4]
  assign _T_259 = 2'h2 == io_reg2dp_y_extension; // @[Mux.scala 46:19:@49.4]
  assign pixel_x_init_w = _T_259 ? _T_252 : {{1'd0}, _T_258}; // @[Mux.scala 46:16:@50.4]
  assign pixel_x_init_offset_w = _T_243 + 6'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 116:80:@52.4]
  assign _T_264 = {pixel_x_stride_w,2'h0}; // @[Cat.scala 30:58:@53.4]
  assign _T_269 = _T_257 ? _T_247 : {{1'd0}, pixel_x_stride_w}; // @[Mux.scala 46:16:@56.4]
  assign pixel_x_add_w = _T_259 ? _T_264 : {{1'd0}, _T_269}; // @[Mux.scala 46:16:@58.4]
  assign pixel_ch_stride_w = {pixel_x_stride_w,6'h0}; // @[Cat.scala 30:58:@59.4]
  assign conv_y_stride_w = io_reg2dp_conv_y_stride_ext + 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 126:74:@60.4]
  assign _T_278 = io_reg2dp_x_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 127:74:@63.4]
  assign x_dilate_w = is_img ? 6'h1 : _T_278; // @[NV_NVDLA_CSC_dl_for_check.scala 127:21:@64.4]
  assign _T_282 = io_reg2dp_y_dilation_ext + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 128:74:@66.4]
  assign y_dilate_w = is_img ? 6'h1 : _T_282; // @[NV_NVDLA_CSC_dl_for_check.scala 128:21:@67.4]
  assign entries_single_w = io_reg2dp_entries + 14'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 144:43:@91.4]
  assign _T_353 = entries_single_w * 15'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 145:41:@93.4]
  assign entries_batch_w = _T_353[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 145:56:@94.4]
  assign entries_w = {{2'd0}, entries_single_w}; // @[NV_NVDLA_CSC_dl_for_check.scala 146:20:@97.4]
  assign h_offset_slice_w = 6'h1 * y_dilate_w; // @[NV_NVDLA_CSC_dl_for_check.scala 147:37:@98.4]
  assign _GEN_684 = {{11'd0}, data_batch}; // @[NV_NVDLA_CSC_dl_for_check.scala 148:33:@99.4]
  assign h_bias_0_stride_w = entries * _GEN_684; // @[NV_NVDLA_CSC_dl_for_check.scala 148:33:@99.4]
  assign _GEN_685 = {{3'd0}, h_offset_slice}; // @[NV_NVDLA_CSC_dl_for_check.scala 149:33:@100.4]
  assign h_bias_1_stride_w = entries * _GEN_685; // @[NV_NVDLA_CSC_dl_for_check.scala 149:33:@100.4]
  assign rls_slices_w = io_reg2dp_rls_slices + 12'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 150:41:@101.4]
  assign _T_360 = io_reg2dp_datain_height_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 151:77:@102.4]
  assign _GEN_686 = {{1'd0}, io_reg2dp_rls_slices}; // @[NV_NVDLA_CSC_dl_for_check.scala 151:113:@103.4]
  assign _T_361 = io_reg2dp_datain_height_ext - _GEN_686; // @[NV_NVDLA_CSC_dl_for_check.scala 151:113:@103.4]
  assign _T_362 = $unsigned(_T_361); // @[NV_NVDLA_CSC_dl_for_check.scala 151:113:@104.4]
  assign slice_left_w = io_reg2dp_skip_data_rls ? _T_360 : _T_362; // @[NV_NVDLA_CSC_dl_for_check.scala 151:23:@105.4]
  assign slices_oprand = layer_st_d1 ? rls_slices : slice_left; // @[NV_NVDLA_CSC_dl_for_check.scala 152:24:@106.4]
  assign _GEN_687 = {{1'd0}, slices_oprand}; // @[NV_NVDLA_CSC_dl_for_check.scala 153:37:@107.4]
  assign slice_entries_w = entries_batch * _GEN_687; // @[NV_NVDLA_CSC_dl_for_check.scala 153:37:@107.4]
  assign _T_547 = is_img ? 34'h3ffffffff : 34'h0; // @[Bitwise.scala 72:12:@178.6]
  assign _T_549 = io_reg2dp_data_bank + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 202:38:@180.6]
  assign _T_554 = io_reg2dp_datain_width_ext + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 203:109:@184.6]
  assign _T_557 = io_reg2dp_weight_channel_ext[12:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 206:109:@190.6]
  assign _T_558 = {{4'd0}, _T_557}; // @[NV_NVDLA_CSC_dl_for_check.scala 206:30:@191.6]
  assign _T_559 = sub_h_total_w[2:1]; // @[NV_NVDLA_CSC_dl_for_check.scala 209:36:@195.6]
  assign _T_562 = {1'h0,io_reg2dp_entries}; // @[Cat.scala 30:58:@224.6]
  assign _GEN_0 = layer_st ? 22'h0 : is_winograd_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_1 = layer_st ? _T_547 : is_img_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_2 = layer_st ? _T_549 : data_bank; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_3 = layer_st ? _T_554 : datain_width; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_4 = layer_st ? io_reg2dp_datain_width_ext : datain_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_5 = layer_st ? io_reg2dp_datain_height_ext : datain_height_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_6 = layer_st ? _T_558 : datain_channel_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_7 = layer_st ? sub_h_total_w : sub_h_total_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_8 = layer_st ? sub_h_total_w : sub_h_total_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_9 = layer_st ? _T_559 : sub_h_total_g2; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_10 = layer_st ? sub_h_total_w : sub_h_total_g3; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_11 = layer_st ? sub_h_total_w : sub_h_total_g4; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_12 = layer_st ? sub_h_total_w : sub_h_total_g5; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_13 = layer_st ? sub_h_total_w : sub_h_total_g6; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_15 = layer_st ? sub_h_total_w : sub_h_total_g8; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_16 = layer_st ? sub_h_total_w : sub_h_total_g9; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_18 = layer_st ? sub_h_total_w : sub_h_total_g11; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_19 = layer_st ? sub_h_cmp_w : sub_h_cmp_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_20 = layer_st ? sub_h_cmp_w : sub_h_cmp_g1; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_21 = layer_st ? conv_x_stride_w : conv_x_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_22 = layer_st ? conv_y_stride_w : conv_y_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_24 = layer_st ? 6'h1 : data_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_25 = layer_st ? 5'h0 : batch_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_26 = layer_st ? pixel_x_init_w : pixel_x_init; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_27 = layer_st ? pixel_x_init_offset_w : pixel_x_init_offset; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_28 = layer_st ? pixel_x_add_w : pixel_x_add; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_29 = layer_st ? {{1'd0}, pixel_x_stride_w} : pixel_x_byte_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_30 = layer_st ? pixel_ch_stride_w : pixel_ch_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_31 = layer_st ? x_dilate_w : x_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_32 = layer_st ? y_dilate_w : y_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_33 = layer_st ? io_reg2dp_pad_value : pad_value; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_34 = layer_st ? entries_w : entries; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_35 = layer_st ? entries_batch_w : entries_batch; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_36 = layer_st ? _T_562 : entries_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_37 = layer_st ? {{2'd0}, h_offset_slice_w} : h_offset_slice; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_38 = layer_st ? {{1'd0}, rls_slices_w} : rls_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_39 = layer_st ? slice_left_w : slice_left; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_40 = layer_st ? io_reg2dp_dataout_width : dataout_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 199:15:@174.4]
  assign _GEN_43 = layer_st_d1 ? h_bias_0_stride_w : h_bias_0_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  assign _GEN_44 = layer_st_d1 ? h_bias_1_stride_w : h_bias_1_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  assign _GEN_45 = layer_st_d1 ? entries : h_bias_2_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  assign _GEN_46 = layer_st_d1 ? entries : h_bias_3_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  assign _GEN_47 = layer_st_d1 ? slice_entries_w : rls_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 244:18:@237.4]
  assign _GEN_48 = is_sg_done ? slice_left : last_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 251:17:@244.4]
  assign _GEN_49 = is_sg_done ? slice_entries_w : last_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 251:17:@244.4]
  assign _T_643 = last_slices != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 315:37:@328.4]
  assign _T_644 = io_sg2dl_reuse_rls & _T_643; // @[NV_NVDLA_CSC_dl_for_check.scala 315:23:@329.4]
  assign _T_1517 = sub_h_total_g3[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 911:32:@1247.4]
  assign _T_1518 = _T_1517 & dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 911:36:@1248.4]
  assign _T_1519 = sub_h_total_g3[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 912:35:@1249.4]
  assign _T_1520 = _T_1519 & dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 912:39:@1250.4]
  assign _T_1521 = _T_1518 | _T_1520; // @[NV_NVDLA_CSC_dl_for_check.scala 911:57:@1251.4]
  assign _T_1522 = sub_h_total_g3[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 913:35:@1252.4]
  assign _T_1523 = _T_1522 & dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 913:39:@1253.4]
  assign dat_rsp_pvld = _T_1521 | _T_1523; // @[NV_NVDLA_CSC_dl_for_check.scala 912:60:@1254.4]
  assign _T_1525 = sub_h_total_g4[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 920:42:@1256.4]
  assign _T_1529 = _T_1525 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1258.4]
  assign _T_1530 = _T_1529 & _T_1507; // @[NV_NVDLA_CSC_dl_for_check.scala 920:47:@1259.4]
  assign _T_1531 = sub_h_total_g4[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 921:42:@1260.4]
  assign _T_1535 = _T_1531 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1262.4]
  assign _T_1536 = _T_1535 & _T_1501; // @[NV_NVDLA_CSC_dl_for_check.scala 921:47:@1263.4]
  assign _T_1537 = _T_1530 | _T_1536; // @[NV_NVDLA_CSC_dl_for_check.scala 920:66:@1264.4]
  assign _T_1538 = sub_h_total_g4[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 922:42:@1265.4]
  assign _T_1542 = _T_1538 ? 27'h7ffffff : 27'h0; // @[Bitwise.scala 72:12:@1267.4]
  assign _T_1543 = _T_1542 & _T_1498; // @[NV_NVDLA_CSC_dl_for_check.scala 922:47:@1268.4]
  assign dat_rsp_pd = _T_1537 | _T_1543; // @[NV_NVDLA_CSC_dl_for_check.scala 921:66:@1269.4]
  assign dat_rsp_rls = dat_rsp_pd[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 946:26:@1288.4]
  assign sub_rls = dat_rsp_pvld & dat_rsp_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 312:29:@327.4]
  assign _T_646 = rls_slices != 14'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 315:66:@330.4]
  assign _T_647 = sub_rls & _T_646; // @[NV_NVDLA_CSC_dl_for_check.scala 315:53:@331.4]
  assign dat_rls = _T_644 | _T_647; // @[NV_NVDLA_CSC_dl_for_check.scala 315:42:@332.4]
  assign sc2cdma_dat_slices_w = sub_rls ? rls_slices : last_slices; // @[NV_NVDLA_CSC_dl_for_check.scala 316:28:@334.4]
  assign _T_650 = sub_rls ? rls_entries : last_entries; // @[NV_NVDLA_CSC_dl_for_check.scala 317:29:@336.4]
  assign sc2cdma_dat_entries_w = _T_650[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 271:34:@266.4 NV_NVDLA_CSC_dl_for_check.scala 317:23:@337.4]
  assign dat_entry_avl_sub = dat_rls ? sc2cdma_dat_entries_w : 15'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 284:28:@278.4]
  assign _T_600 = dat_entry_st + dat_entry_avl_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 289:37:@283.4]
  assign dat_entry_st_inc = dat_entry_st + dat_entry_avl_sub; // @[NV_NVDLA_CSC_dl_for_check.scala 289:37:@284.4]
  assign _T_606 = {data_bank,9'h0}; // @[Cat.scala 30:58:@286.4]
  assign _T_607 = dat_entry_st_inc - _T_606; // @[NV_NVDLA_CSC_dl_for_check.scala 290:46:@287.4]
  assign _T_608 = $unsigned(_T_607); // @[NV_NVDLA_CSC_dl_for_check.scala 290:46:@288.4]
  assign dat_entry_st_inc_wrap = _T_608[14:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 290:46:@289.4]
  assign is_dat_entry_st_wrap = dat_entry_st_inc >= _T_606; // @[NV_NVDLA_CSC_dl_for_check.scala 291:45:@292.4]
  assign _T_616 = is_dat_entry_st_wrap ? dat_entry_st_inc_wrap : dat_entry_st_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 292:83:@293.4]
  assign dat_entry_st_w = io_sc2cdma_dat_pending_req ? 15'h0 : _T_616; // @[NV_NVDLA_CSC_dl_for_check.scala 292:25:@294.4]
  assign _T_638 = dat_rls | io_sc2cdma_dat_pending_req; // @[NV_NVDLA_CSC_dl_for_check.scala 303:13:@317.4]
  assign _GEN_55 = _T_638 ? dat_entry_st_w : dat_entry_st; // @[NV_NVDLA_CSC_dl_for_check.scala 303:25:@318.4]
  assign _GEN_57 = dat_rls ? sc2cdma_dat_slices_w : _T_656; // @[Reg.scala 20:19:@342.4]
  assign _GEN_58 = dat_rls ? sc2cdma_dat_entries_w : _T_659; // @[Reg.scala 20:19:@347.4]
  assign _GEN_59 = io_sg2dl_pd_valid ? io_sg2dl_pd_bits : _T_681; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@366.4]
  assign _GEN_60 = _T_664 ? _T_681 : _T_684; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@370.4]
  assign _GEN_61 = _T_667 ? _T_684 : _T_687; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@374.4]
  assign _GEN_62 = _T_670 ? _T_687 : _T_690; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@378.4]
  assign _GEN_63 = _T_673 ? _T_690 : _T_693; // @[NV_NVDLA_CSC_dl_for_check.scala 342:26:@382.4]
  assign _T_694 = is_winograd_d1[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 347:36:@385.4]
  assign dl_in_pvld = _T_694 ? io_sg2dl_pd_valid : _T_676; // @[NV_NVDLA_CSC_dl_for_check.scala 347:21:@386.4]
  assign _T_695 = is_winograd_d1[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 348:34:@387.4]
  assign dl_in_pd = _T_695 ? io_sg2dl_pd_bits : _T_693; // @[NV_NVDLA_CSC_dl_for_check.scala 348:19:@388.4]
  assign _GEN_64 = dl_in_pvld ? dl_in_pd : _T_714; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@402.4]
  assign _GEN_65 = _T_700 ? _T_714 : _T_717; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@406.4]
  assign _GEN_66 = _T_703 ? _T_717 : _T_720; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@410.4]
  assign _GEN_67 = _T_706 ? _T_720 : _T_723; // @[NV_NVDLA_CSC_dl_for_check.scala 361:23:@414.4]
  assign _T_724 = sub_h_total_g0[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 366:30:@417.4]
  assign _T_725 = _T_724 & _T_700; // @[NV_NVDLA_CSC_dl_for_check.scala 366:34:@418.4]
  assign _T_726 = sub_h_total_g0[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 367:30:@419.4]
  assign _T_727 = _T_726 & _T_706; // @[NV_NVDLA_CSC_dl_for_check.scala 367:34:@420.4]
  assign _T_728 = _T_725 | _T_727; // @[NV_NVDLA_CSC_dl_for_check.scala 366:50:@421.4]
  assign _T_729 = sub_h_total_g0[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 368:30:@422.4]
  assign _T_730 = _T_729 & _T_709; // @[NV_NVDLA_CSC_dl_for_check.scala 368:34:@423.4]
  assign dl_pvld = _T_728 | _T_730; // @[NV_NVDLA_CSC_dl_for_check.scala 367:50:@424.4]
  assign _T_731 = sub_h_total_g1[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 370:37:@425.4]
  assign _T_735 = _T_731 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@427.4]
  assign _T_736 = _T_735 & _T_714; // @[NV_NVDLA_CSC_dl_for_check.scala 370:42:@428.4]
  assign _T_737 = sub_h_total_g1[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 371:37:@429.4]
  assign _T_741 = _T_737 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@431.4]
  assign _T_742 = _T_741 & _T_720; // @[NV_NVDLA_CSC_dl_for_check.scala 371:42:@432.4]
  assign _T_743 = _T_736 | _T_742; // @[NV_NVDLA_CSC_dl_for_check.scala 370:56:@433.4]
  assign _T_744 = sub_h_total_g1[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 372:37:@434.4]
  assign _T_748 = _T_744 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12:@436.4]
  assign _T_749 = _T_748 & _T_723; // @[NV_NVDLA_CSC_dl_for_check.scala 372:42:@437.4]
  assign dl_pd = _T_743 | _T_749; // @[NV_NVDLA_CSC_dl_for_check.scala 371:56:@438.4]
  assign dl_w_offset = dl_pd[4:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 375:24:@439.4]
  assign dl_h_offset = dl_pd[9:5]; // @[NV_NVDLA_CSC_dl_for_check.scala 376:24:@440.4]
  assign dl_channel_size = dl_pd[16:10]; // @[NV_NVDLA_CSC_dl_for_check.scala 377:28:@441.4]
  assign dl_stripe_length = dl_pd[23:17]; // @[NV_NVDLA_CSC_dl_for_check.scala 378:29:@442.4]
  assign dl_cur_sub_h = dl_pd[25:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 379:25:@443.4]
  assign dl_block_end = dl_pd[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 380:25:@444.4]
  assign dl_channel_end = dl_pd[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 381:27:@445.4]
  assign dl_group_end = dl_pd[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 382:25:@446.4]
  assign dl_layer_end = dl_pd[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 383:25:@447.4]
  assign dl_dat_release = dl_pd[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 384:27:@448.4]
  assign _T_806 = stripe_cnt != 7'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 439:37:@505.4]
  assign _T_807 = ~ _T_806; // @[NV_NVDLA_CSC_dl_for_check.scala 439:24:@506.4]
  assign _T_809 = sub_h_cnt != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 439:56:@507.4]
  assign _T_810 = ~ _T_809; // @[NV_NVDLA_CSC_dl_for_check.scala 439:44:@508.4]
  assign _T_811 = _T_807 & _T_810; // @[NV_NVDLA_CSC_dl_for_check.scala 439:42:@509.4]
  assign _T_813 = batch_cnt != 5'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 439:75:@510.4]
  assign _T_814 = ~ _T_813; // @[NV_NVDLA_CSC_dl_for_check.scala 439:63:@511.4]
  assign _T_815 = _T_811 & _T_814; // @[NV_NVDLA_CSC_dl_for_check.scala 439:61:@512.4]
  assign _T_817 = _T_815 ? 1'h0 : dat_exec_valid_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 439:22:@513.4]
  assign dat_exec_valid = dl_pvld ? 1'h1 : _T_817; // @[NV_NVDLA_CSC_dl_for_check.scala 438:22:@514.4]
  assign _T_754 = layer_st | dat_exec_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 391:15:@452.4]
  assign _T_758 = batch_cnt + 5'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 394:28:@454.6]
  assign is_batch_end = batch_cnt == batch_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 398:27:@459.4]
  assign _T_759 = is_batch_end ? 6'h0 : _T_758; // @[NV_NVDLA_CSC_dl_for_check.scala 393:21:@455.6]
  assign _T_760 = layer_st ? 6'h0 : _T_759; // @[NV_NVDLA_CSC_dl_for_check.scala 392:21:@456.6]
  assign _GEN_68 = _T_754 ? _T_760 : {{1'd0}, batch_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 391:32:@453.4]
  assign sub_h_cnt_inc = sub_h_cnt + 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 404:31:@463.4]
  assign is_sub_h_end = sub_h_cnt_inc == sub_h_cmp_g0; // @[NV_NVDLA_CSC_dl_for_check.scala 405:32:@464.4]
  assign _T_767 = is_winograd_d1[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 406:51:@466.4]
  assign _T_769 = io_reg2dp_y_extension != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 406:82:@467.4]
  assign _T_770 = _T_767 | _T_769; // @[NV_NVDLA_CSC_dl_for_check.scala 406:55:@468.4]
  assign _T_771 = _T_770 & dat_exec_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 406:88:@469.4]
  assign sub_h_cnt_reg_en = layer_st | _T_771; // @[NV_NVDLA_CSC_dl_for_check.scala 406:33:@470.4]
  assign _T_772 = layer_st | is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 408:31:@472.6]
  assign _T_774 = _T_772 ? 3'h0 : sub_h_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 408:21:@473.6]
  assign _GEN_69 = sub_h_cnt_reg_en ? _T_774 : {{1'd0}, sub_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 407:23:@471.4]
  assign _T_780 = stripe_cnt + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 416:34:@479.4]
  assign stripe_cnt_inc = _T_780[6:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 416:41:@480.4]
  assign _T_781 = stripe_cnt_inc == dl_stripe_length; // @[NV_NVDLA_CSC_dl_for_check.scala 417:51:@481.4]
  assign is_stripe_equal = is_batch_end & _T_781; // @[NV_NVDLA_CSC_dl_for_check.scala 417:33:@482.4]
  assign is_stripe_end = is_stripe_equal & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 418:34:@484.4]
  assign _T_784 = dat_exec_valid & is_batch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 419:52:@486.4]
  assign stripe_cnt_reg_en = layer_st | _T_784; // @[NV_NVDLA_CSC_dl_for_check.scala 419:34:@487.4]
  assign _T_786 = ~ is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 423:41:@489.6]
  assign _T_787 = is_stripe_equal & _T_786; // @[NV_NVDLA_CSC_dl_for_check.scala 423:39:@490.6]
  assign _T_789 = is_stripe_end ? 7'h0 : stripe_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 424:22:@491.6]
  assign _T_790 = _T_787 ? stripe_cnt : _T_789; // @[NV_NVDLA_CSC_dl_for_check.scala 423:22:@492.6]
  assign _T_791 = layer_st ? 7'h0 : _T_790; // @[NV_NVDLA_CSC_dl_for_check.scala 422:22:@493.6]
  assign _GEN_70 = stripe_cnt_reg_en ? _T_791 : stripe_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 421:24:@488.4]
  assign dat_pipe_valid = dl_pvld | dat_pipe_local_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 437:27:@503.4]
  assign _T_799 = dat_pipe_valid & is_stripe_equal; // @[NV_NVDLA_CSC_dl_for_check.scala 434:49:@500.4]
  assign _T_802 = dl_pvld ? 1'h1 : dat_pipe_local_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 435:32:@501.4]
  assign dat_pipe_local_valid_w = _T_799 ? 1'h0 : _T_802; // @[NV_NVDLA_CSC_dl_for_check.scala 434:33:@502.4]
  assign dat_req_bytes = {1'h0,dl_channel_size}; // @[Cat.scala 30:58:@520.4]
  assign _GEN_71 = dat_exec_valid ? dat_req_bytes : dat_req_bytes_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 449:21:@521.4]
  assign _GEN_690 = {{10'd0}, sub_h_cmp_g1}; // @[NV_NVDLA_CSC_dl_for_check.scala 459:39:@526.4]
  assign _T_826 = dataout_w_cnt + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 459:39:@526.4]
  assign dataout_w_cnt_inc = dataout_w_cnt + _GEN_690; // @[NV_NVDLA_CSC_dl_for_check.scala 459:39:@527.4]
  assign _T_827 = is_batch_end & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 460:29:@528.4]
  assign _T_828 = dataout_w_cnt >= dataout_width_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 460:61:@529.4]
  assign is_w_end = _T_827 & _T_828; // @[NV_NVDLA_CSC_dl_for_check.scala 460:44:@530.4]
  assign _T_830 = ~ dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 463:43:@533.4]
  assign _T_831 = is_stripe_end & _T_830; // @[NV_NVDLA_CSC_dl_for_check.scala 463:41:@534.4]
  assign _T_832 = is_w_end ? {{9'd0}, dataout_w_init} : dataout_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 464:26:@535.4]
  assign _T_833 = _T_831 ? dataout_w_ori : _T_832; // @[NV_NVDLA_CSC_dl_for_check.scala 463:26:@536.4]
  assign dataout_w_cnt_w = layer_st ? {{9'd0}, dataout_w_init} : _T_833; // @[NV_NVDLA_CSC_dl_for_check.scala 462:26:@537.4]
  assign _T_835 = _T_784 & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 465:70:@539.4]
  assign dataout_w_cnt_reg_en = layer_st | _T_835; // @[NV_NVDLA_CSC_dl_for_check.scala 465:37:@540.4]
  assign _T_836 = dat_exec_valid & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 466:55:@541.4]
  assign _T_837 = _T_836 & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 466:71:@542.4]
  assign dataout_w_ori_reg_en = layer_st | _T_837; // @[NV_NVDLA_CSC_dl_for_check.scala 466:37:@543.4]
  assign _GEN_72 = dataout_w_cnt_reg_en ? dataout_w_cnt_w : dataout_w_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 468:27:@544.4]
  assign _GEN_73 = dataout_w_ori_reg_en ? dataout_w_cnt_w : dataout_w_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 471:27:@547.4]
  assign is_last_channel = datain_c_cnt == datain_channel_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 478:37:@551.4]
  assign _T_841 = _T_836 & dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 479:70:@553.4]
  assign datain_c_cnt_reg_en = layer_st | _T_841; // @[NV_NVDLA_CSC_dl_for_check.scala 479:36:@554.4]
  assign _T_845 = datain_c_cnt + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 484:34:@556.6]
  assign _T_846 = datain_c_cnt + 11'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 484:34:@557.6]
  assign _T_847 = dl_channel_end ? 11'h0 : _T_846; // @[NV_NVDLA_CSC_dl_for_check.scala 483:24:@558.6]
  assign _T_848 = layer_st ? 11'h0 : _T_847; // @[NV_NVDLA_CSC_dl_for_check.scala 482:24:@559.6]
  assign _GEN_74 = datain_c_cnt_reg_en ? _T_848 : datain_c_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 481:26:@555.4]
  assign _GEN_691 = {{8'd0}, io_reg2dp_pad_left}; // @[NV_NVDLA_CSC_dl_for_check.scala 500:41:@571.4]
  assign _T_869 = 13'h0 - _GEN_691; // @[NV_NVDLA_CSC_dl_for_check.scala 500:41:@571.4]
  assign _T_870 = $unsigned(_T_869); // @[NV_NVDLA_CSC_dl_for_check.scala 500:41:@572.4]
  assign datain_w_cnt_st = is_img ? 14'h0 : _T_870; // @[NV_NVDLA_CSC_dl_for_check.scala 498:26:@574.4]
  assign _T_872 = is_winograd_d1[3]; // @[NV_NVDLA_CSC_dl_for_check.scala 501:42:@575.4]
  assign _T_874 = datain_w_cnt + 14'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 501:60:@576.4]
  assign _GEN_692 = {{10'd0}, conv_x_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 501:81:@577.4]
  assign _T_875 = datain_w_cnt + _GEN_692; // @[NV_NVDLA_CSC_dl_for_check.scala 501:81:@577.4]
  assign datain_w_cnt_inc = _T_872 ? _T_874 : _T_875; // @[NV_NVDLA_CSC_dl_for_check.scala 501:27:@578.4]
  assign _T_878 = is_w_end ? {{1'd0}, datain_w_cnt_st} : datain_w_cnt_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 506:25:@581.4]
  assign _T_879 = _T_831 ? {{1'd0}, datain_w_ori} : _T_878; // @[NV_NVDLA_CSC_dl_for_check.scala 505:25:@582.4]
  assign datain_w_cnt_w = layer_st ? {{1'd0}, datain_w_cnt_st} : _T_879; // @[NV_NVDLA_CSC_dl_for_check.scala 504:25:@583.4]
  assign _GEN_693 = {{1'd0}, dl_w_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 508:35:@584.4]
  assign dl_w_offset_ext = _GEN_693 * x_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 508:35:@584.4]
  assign _GEN_694 = {{3'd0}, dl_w_offset_ext}; // @[NV_NVDLA_CSC_dl_for_check.scala 509:34:@585.4]
  assign _T_880 = datain_w_cnt + _GEN_694; // @[NV_NVDLA_CSC_dl_for_check.scala 509:34:@585.4]
  assign datain_w_cur = _T_880[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 509:53:@586.4]
  assign _T_883 = is_img_d1[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 510:96:@589.4]
  assign _T_884 = ~ _T_883; // @[NV_NVDLA_CSC_dl_for_check.scala 510:86:@590.4]
  assign _T_885 = _T_835 & _T_884; // @[NV_NVDLA_CSC_dl_for_check.scala 510:84:@591.4]
  assign datain_w_cnt_reg_en = layer_st | _T_885; // @[NV_NVDLA_CSC_dl_for_check.scala 510:36:@592.4]
  assign _T_888 = is_img_d1[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 511:99:@595.4]
  assign _T_889 = ~ _T_888; // @[NV_NVDLA_CSC_dl_for_check.scala 511:89:@596.4]
  assign _T_890 = _T_837 & _T_889; // @[NV_NVDLA_CSC_dl_for_check.scala 511:87:@597.4]
  assign datain_w_ori_reg_en = layer_st | _T_890; // @[NV_NVDLA_CSC_dl_for_check.scala 511:36:@598.4]
  assign pixel_x_cnt_add = is_sub_h_end ? pixel_x_add : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 514:26:@599.4]
  assign _T_894 = _T_243 == 6'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 516:79:@601.4]
  assign _T_898 = _T_557 + 7'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 517:75:@604.4]
  assign total_channel_op = _T_894 ? {{1'd0}, _T_557} : _T_898; // @[NV_NVDLA_CSC_dl_for_check.scala 516:27:@605.4]
  assign _T_899 = dl_channel_end & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 518:37:@606.4]
  assign _T_901 = dl_block_end & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 519:35:@607.4]
  assign _T_903 = channel_op_cnt + 13'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 519:66:@608.4]
  assign _T_904 = _T_901 ? _T_903 : {{1'd0}, channel_op_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 519:22:@609.4]
  assign _T_905 = _T_899 ? 14'h2 : _T_904; // @[NV_NVDLA_CSC_dl_for_check.scala 518:22:@610.4]
  assign _GEN_695 = {{5'd0}, total_channel_op}; // @[NV_NVDLA_CSC_dl_for_check.scala 521:44:@612.4]
  assign next_is_last_channel = channel_op_cnt >= _GEN_695; // @[NV_NVDLA_CSC_dl_for_check.scala 521:44:@612.4]
  assign _T_906 = is_stripe_end & dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 525:39:@613.4]
  assign _T_907 = _T_906 & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 525:54:@614.4]
  assign _T_908 = _T_907 & is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 525:71:@615.4]
  assign _T_911 = ~ is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 526:73:@618.4]
  assign _T_912 = _T_907 & _T_911; // @[NV_NVDLA_CSC_dl_for_check.scala 526:71:@619.4]
  assign _GEN_696 = {{4'd0}, pixel_ch_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 526:99:@620.4]
  assign _T_913 = pixel_w_ch_ori + _GEN_696; // @[NV_NVDLA_CSC_dl_for_check.scala 526:99:@620.4]
  assign _T_915 = _T_906 & next_is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 527:54:@622.4]
  assign _GEN_697 = {{9'd0}, pixel_x_init_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 527:90:@623.4]
  assign _T_916 = pixel_w_ori + _GEN_697; // @[NV_NVDLA_CSC_dl_for_check.scala 527:90:@623.4]
  assign _T_918 = ~ next_is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 528:56:@625.4]
  assign _T_919 = _T_906 & _T_918; // @[NV_NVDLA_CSC_dl_for_check.scala 528:54:@626.4]
  assign _T_921 = pixel_w_ori + 16'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 528:91:@627.4]
  assign _T_922 = ~ dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 529:41:@628.4]
  assign _T_923 = is_stripe_end & _T_922; // @[NV_NVDLA_CSC_dl_for_check.scala 529:39:@629.4]
  assign _GEN_698 = {{8'd0}, pixel_x_cnt_add}; // @[NV_NVDLA_CSC_dl_for_check.scala 529:81:@630.4]
  assign _T_924 = pixel_w_cnt + _GEN_698; // @[NV_NVDLA_CSC_dl_for_check.scala 529:81:@630.4]
  assign _T_925 = _T_923 ? {{1'd0}, pixel_w_ori} : _T_924; // @[NV_NVDLA_CSC_dl_for_check.scala 529:24:@631.4]
  assign _T_926 = _T_919 ? _T_921 : _T_925; // @[NV_NVDLA_CSC_dl_for_check.scala 528:24:@632.4]
  assign _T_927 = _T_915 ? _T_916 : _T_926; // @[NV_NVDLA_CSC_dl_for_check.scala 527:24:@633.4]
  assign _T_928 = _T_912 ? _T_913 : _T_927; // @[NV_NVDLA_CSC_dl_for_check.scala 526:24:@634.4]
  assign _T_929 = _T_908 ? {{10'd0}, pixel_x_init} : _T_928; // @[NV_NVDLA_CSC_dl_for_check.scala 525:24:@635.4]
  assign pixel_w_cnt_w = layer_st_d1 ? {{10'd0}, pixel_x_init} : _T_929; // @[NV_NVDLA_CSC_dl_for_check.scala 524:24:@636.4]
  assign _T_935 = pixel_w_cnt[15:6]; // @[NV_NVDLA_CSC_dl_for_check.scala 531:68:@638.4]
  assign pixel_w_cur = {5'h0,_T_935}; // @[Cat.scala 30:58:@639.4]
  assign _T_944 = is_img_d1[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 534:68:@650.4]
  assign _T_945 = dat_exec_valid & _T_944; // @[NV_NVDLA_CSC_dl_for_check.scala 534:57:@651.4]
  assign _T_946 = _T_945 & is_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 534:72:@652.4]
  assign _T_947 = _T_946 & dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 534:88:@653.4]
  assign _T_948 = _T_947 & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 534:103:@654.4]
  assign pixel_ch_ori_reg_en = layer_st_d1 | _T_948; // @[NV_NVDLA_CSC_dl_for_check.scala 534:39:@655.4]
  assign _T_950 = _T_883 & dl_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 536:42:@657.4]
  assign _T_953 = pixel_force_clr_d1 ? 1'h0 : pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 536:74:@658.4]
  assign pixel_force_fetch = _T_950 ? 1'h1 : _T_953; // @[NV_NVDLA_CSC_dl_for_check.scala 536:28:@659.4]
  assign _T_955 = _T_883 & is_sub_h_end; // @[NV_NVDLA_CSC_dl_for_check.scala 537:36:@661.4]
  assign _T_956 = pixel_force_fetch | pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 537:72:@662.4]
  assign pixel_force_clr = _T_955 & _T_956; // @[NV_NVDLA_CSC_dl_for_check.scala 537:51:@663.4]
  assign _GEN_75 = datain_w_cnt_reg_en ? datain_w_cnt_w : {{1'd0}, datain_w_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 539:26:@664.4]
  assign _GEN_76 = datain_w_cnt_reg_en ? pixel_w_cnt_w : {{1'd0}, pixel_w_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 539:26:@664.4]
  assign _GEN_77 = datain_w_ori_reg_en ? datain_w_cnt_w : {{1'd0}, datain_w_ori}; // @[NV_NVDLA_CSC_dl_for_check.scala 543:26:@668.4]
  assign _GEN_78 = datain_w_ori_reg_en ? pixel_w_cnt_w : {{1'd0}, pixel_w_ori}; // @[NV_NVDLA_CSC_dl_for_check.scala 543:26:@668.4]
  assign _GEN_79 = pixel_ch_ori_reg_en ? pixel_w_cnt_w : {{1'd0}, pixel_w_ch_ori}; // @[NV_NVDLA_CSC_dl_for_check.scala 547:26:@672.4]
  assign _GEN_699 = {{9'd0}, io_reg2dp_pad_top}; // @[NV_NVDLA_CSC_dl_for_check.scala 556:77:@677.4]
  assign _T_963 = 14'h0 - _GEN_699; // @[NV_NVDLA_CSC_dl_for_check.scala 556:77:@677.4]
  assign datain_h_cnt_st = $unsigned(_T_963); // @[NV_NVDLA_CSC_dl_for_check.scala 556:77:@678.4]
  assign _GEN_700 = {{10'd0}, conv_y_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 557:37:@680.4]
  assign _T_965 = datain_h_cnt + _GEN_700; // @[NV_NVDLA_CSC_dl_for_check.scala 557:37:@680.4]
  assign datain_h_cnt_inc = datain_h_cnt + _GEN_700; // @[NV_NVDLA_CSC_dl_for_check.scala 557:37:@681.4]
  assign _T_966 = is_stripe_end & dl_group_end; // @[NV_NVDLA_CSC_dl_for_check.scala 558:52:@682.4]
  assign _T_967 = layer_st | _T_966; // @[NV_NVDLA_CSC_dl_for_check.scala 558:35:@683.4]
  assign _T_970 = is_w_end ? datain_h_cnt_inc : datain_h_cnt; // @[NV_NVDLA_CSC_dl_for_check.scala 560:25:@686.4]
  assign _T_971 = _T_831 ? datain_h_ori : _T_970; // @[NV_NVDLA_CSC_dl_for_check.scala 559:25:@687.4]
  assign datain_h_cnt_w = _T_967 ? datain_h_cnt_st : {{1'd0}, _T_971}; // @[NV_NVDLA_CSC_dl_for_check.scala 558:25:@688.4]
  assign _T_974 = _T_831 | is_w_end; // @[NV_NVDLA_CSC_dl_for_check.scala 561:91:@691.4]
  assign _T_975 = dat_exec_valid & _T_974; // @[NV_NVDLA_CSC_dl_for_check.scala 561:54:@692.4]
  assign datain_h_cnt_reg_en = layer_st | _T_975; // @[NV_NVDLA_CSC_dl_for_check.scala 561:36:@693.4]
  assign _GEN_701 = {{1'd0}, dl_h_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 563:35:@697.4]
  assign dl_h_offset_ext = _GEN_701 * y_dilate; // @[NV_NVDLA_CSC_dl_for_check.scala 563:35:@697.4]
  assign _GEN_702 = {{3'd0}, dl_h_offset_ext}; // @[NV_NVDLA_CSC_dl_for_check.scala 564:34:@698.4]
  assign _T_978 = datain_h_cnt + _GEN_702; // @[NV_NVDLA_CSC_dl_for_check.scala 564:34:@698.4]
  assign _GEN_703 = {{13'd0}, sub_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 564:53:@699.4]
  assign _T_979 = _T_978 + _GEN_703; // @[NV_NVDLA_CSC_dl_for_check.scala 564:53:@699.4]
  assign datain_h_cur = _T_979[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 564:66:@700.4]
  assign _GEN_80 = datain_h_cnt_reg_en ? datain_h_cnt_w : {{1'd0}, datain_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 566:26:@701.4]
  assign _GEN_81 = dataout_w_ori_reg_en ? datain_h_cnt_w : {{1'd0}, datain_h_ori}; // @[NV_NVDLA_CSC_dl_for_check.scala 567:26:@704.4]
  assign _T_980 = datain_w_cur[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 570:39:@707.4]
  assign _GEN_704 = {{1'd0}, datain_width_cmp}; // @[NV_NVDLA_CSC_dl_for_check.scala 570:59:@708.4]
  assign _T_981 = datain_w_cur > _GEN_704; // @[NV_NVDLA_CSC_dl_for_check.scala 570:59:@708.4]
  assign _T_982 = _T_980 | _T_981; // @[NV_NVDLA_CSC_dl_for_check.scala 570:44:@709.4]
  assign _T_983 = datain_h_cur[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 570:92:@710.4]
  assign _T_984 = _T_982 | _T_983; // @[NV_NVDLA_CSC_dl_for_check.scala 570:78:@711.4]
  assign _GEN_705 = {{1'd0}, datain_height_cmp}; // @[NV_NVDLA_CSC_dl_for_check.scala 570:112:@712.4]
  assign _T_985 = datain_h_cur > _GEN_705; // @[NV_NVDLA_CSC_dl_for_check.scala 570:112:@712.4]
  assign dat_conv_req_dummy = _T_984 | _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 570:97:@713.4]
  assign _T_986 = datain_w_cur[13:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 572:35:@714.4]
  assign _T_988 = _T_986 != 12'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 572:43:@715.4]
  assign _T_989 = datain_w_cur[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 572:61:@716.4]
  assign _T_990 = _T_988 & _T_989; // @[NV_NVDLA_CSC_dl_for_check.scala 572:47:@717.4]
  assign _T_991 = stripe_cnt[6:1]; // @[NV_NVDLA_CSC_dl_for_check.scala 572:77:@718.4]
  assign _T_993 = _T_991 != 6'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 572:84:@719.4]
  assign dat_wg_req_skip = _T_990 & _T_993; // @[NV_NVDLA_CSC_dl_for_check.scala 572:65:@720.4]
  assign dat_img_req_dummy = _T_983 | _T_985; // @[NV_NVDLA_CSC_dl_for_check.scala 573:42:@723.4]
  assign _T_1080 = is_img_d1[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 659:33:@821.4]
  assign _T_1081 = is_winograd_d1[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 660:38:@822.4]
  assign _T_1082 = ~ is_last_channel; // @[NV_NVDLA_CSC_dl_for_check.scala 661:24:@823.4]
  assign _T_1084 = _T_1082 | _T_1081; // @[NV_NVDLA_CSC_dl_for_check.scala 661:41:@825.4]
  assign _T_1086 = datain_w_cur[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 661:97:@826.4]
  assign _T_1087 = {2'h0,_T_1086}; // @[Cat.scala 30:58:@827.4]
  assign _T_1089 = dat_req_bytes > 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 662:38:@828.4]
  assign _T_1094 = datain_w_cur[12:1]; // @[NV_NVDLA_CSC_dl_for_check.scala 663:54:@831.4]
  assign _T_1095 = {3'h0,_T_1094}; // @[Cat.scala 30:58:@832.4]
  assign _T_1096 = _T_1089 ? _T_1087 : _T_1095; // @[NV_NVDLA_CSC_dl_for_check.scala 662:23:@833.4]
  assign _T_1097 = _T_1084 ? _T_1087 : _T_1096; // @[NV_NVDLA_CSC_dl_for_check.scala 661:23:@834.4]
  assign _T_1098 = _T_1081 ? {{1'd0}, datain_w_cnt} : _T_1097; // @[NV_NVDLA_CSC_dl_for_check.scala 660:23:@835.4]
  assign w_bias_int8 = _T_1080 ? pixel_w_cur : _T_1098; // @[NV_NVDLA_CSC_dl_for_check.scala 659:23:@836.4]
  assign w_bias_w = w_bias_int8[13:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 673:24:@838.4]
  assign _T_997 = w_bias_w[13:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 577:32:@725.4]
  assign _GEN_707 = {{3'd0}, _T_997}; // @[NV_NVDLA_CSC_dl_for_check.scala 577:40:@726.4]
  assign dat_img_req_skip = _GEN_707 > entries_cmp; // @[NV_NVDLA_CSC_dl_for_check.scala 577:40:@726.4]
  assign _T_998 = is_img_d1[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 578:34:@727.4]
  assign _T_999 = is_winograd_d1[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 578:76:@728.4]
  assign _T_1000 = _T_999 ? 1'h0 : dat_conv_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 578:61:@729.4]
  assign dat_req_dummy = _T_998 ? dat_img_req_dummy : _T_1000; // @[NV_NVDLA_CSC_dl_for_check.scala 578:24:@730.4]
  assign _T_1001 = is_winograd_d1[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 579:35:@731.4]
  assign _T_1002 = _T_1001 & dat_wg_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 579:39:@732.4]
  assign _T_1003 = is_img_d1[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 579:70:@733.4]
  assign _T_1004 = _T_1003 & dat_img_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 579:74:@734.4]
  assign dat_req_skip = _T_1002 | _T_1004; // @[NV_NVDLA_CSC_dl_for_check.scala 579:58:@735.4]
  assign _T_1005 = ~ dat_req_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 580:39:@736.4]
  assign _T_1006 = dat_exec_valid & _T_1005; // @[NV_NVDLA_CSC_dl_for_check.scala 580:37:@737.4]
  assign _T_1007 = ~ dat_req_skip; // @[NV_NVDLA_CSC_dl_for_check.scala 580:56:@738.4]
  assign dat_req_valid = _T_1006 & _T_1007; // @[NV_NVDLA_CSC_dl_for_check.scala 580:54:@739.4]
  assign _T_1008 = is_img_d1[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 583:37:@740.4]
  assign _T_1009 = ~ _T_1008; // @[NV_NVDLA_CSC_dl_for_check.scala 583:27:@741.4]
  assign _T_1010 = datain_c_cnt[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 583:54:@742.4]
  assign dat_req_sub_c_w = _T_1009 ? _T_1010 : dl_block_end; // @[NV_NVDLA_CSC_dl_for_check.scala 583:26:@743.4]
  assign _T_1011 = is_winograd_d1[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 584:41:@744.4]
  assign _T_1013 = ~ _T_989; // @[NV_NVDLA_CSC_dl_for_check.scala 584:46:@746.4]
  assign _T_1014 = datain_w_cur[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 584:76:@747.4]
  assign dat_req_sub_w_w = _T_1011 ? {{1'd0}, _T_1013} : _T_1014; // @[NV_NVDLA_CSC_dl_for_check.scala 584:26:@748.4]
  assign _T_1016 = sub_h_cnt == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 585:55:@749.4]
  assign dat_req_sub_w_st_en = dat_exec_valid & _T_1016; // @[NV_NVDLA_CSC_dl_for_check.scala 585:42:@750.4]
  assign dat_req_stripe_end = is_stripe_equal & dat_pipe_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 588:42:@752.4]
  assign dat_req_flag_w = {dl_layer_end,dl_channel_end,dat_req_stripe_end,dl_pvld,batch_cnt}; // @[Cat.scala 30:58:@756.4]
  assign _T_1040 = dl_dat_release & is_stripe_equal; // @[NV_NVDLA_CSC_dl_for_check.scala 615:38:@776.6]
  assign _T_1041 = _T_1040 & dat_pipe_valid; // @[NV_NVDLA_CSC_dl_for_check.scala 615:56:@777.6]
  assign _GEN_82 = dat_exec_valid ? dat_req_sub_w_w : dat_req_sub_w_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_83 = dat_exec_valid ? sub_h_cnt : dat_req_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_84 = dat_exec_valid ? dat_req_sub_c_w : dat_req_sub_c_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_85 = dat_exec_valid ? is_last_channel : dat_req_ch_end_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_86 = dat_exec_valid ? dat_req_dummy : dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_87 = dat_exec_valid ? dl_cur_sub_h : dat_req_cur_sub_h_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_88 = dat_exec_valid ? dat_req_flag_w : dat_req_flag_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_89 = dat_exec_valid ? _T_1041 : dat_req_rls_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_90 = dat_exec_valid ? pixel_force_fetch : pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_91 = dat_exec_valid ? pixel_force_clr : pixel_force_clr_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 607:21:@768.4]
  assign _GEN_92 = dat_req_sub_w_st_en ? dl_pvld : dat_req_sub_w_st_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 619:26:@782.4]
  assign _T_1056 = is_img_d1[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 636:32:@792.4]
  assign _T_1057 = ~ _T_1056; // @[NV_NVDLA_CSC_dl_for_check.scala 636:22:@793.4]
  assign _T_1058 = datain_width[11:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 636:49:@794.4]
  assign c_bias_add = _T_1057 ? _T_1058 : 12'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 636:21:@795.4]
  assign _T_1061 = is_stripe_end & dl_channel_end; // @[NV_NVDLA_CSC_dl_for_check.scala 638:34:@796.4]
  assign _GEN_708 = {{1'd0}, c_bias_add}; // @[NV_NVDLA_CSC_dl_for_check.scala 638:64:@797.4]
  assign _T_1063 = c_bias + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 638:64:@797.4]
  assign _T_1064 = c_bias + _GEN_708; // @[NV_NVDLA_CSC_dl_for_check.scala 638:64:@798.4]
  assign _T_1065 = _T_1061 ? 13'h0 : _T_1064; // @[NV_NVDLA_CSC_dl_for_check.scala 638:19:@799.4]
  assign c_bias_w = layer_st ? 13'h0 : _T_1065; // @[NV_NVDLA_CSC_dl_for_check.scala 637:19:@800.4]
  assign c_bias_d1_reg_en = c_bias != c_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 640:31:@804.4]
  assign _GEN_709 = {{9'd0}, datain_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 643:32:@805.4]
  assign _T_1068 = _GEN_709 * h_bias_0_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 643:32:@805.4]
  assign h_bias_0_w = _T_1068[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 643:50:@806.4]
  assign _GEN_710 = {{26'd0}, dl_h_offset}; // @[NV_NVDLA_CSC_dl_for_check.scala 644:31:@807.4]
  assign _T_1069 = _GEN_710 * h_bias_1_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 644:31:@807.4]
  assign h_bias_1_w = _T_1069[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 644:49:@808.4]
  assign _GEN_711 = {{12'd0}, batch_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 645:29:@809.4]
  assign _T_1070 = _GEN_711 * h_bias_2_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 645:29:@809.4]
  assign h_bias_2_w = _T_1070[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 645:47:@810.4]
  assign _GEN_712 = {{15'd0}, sub_h_cnt}; // @[NV_NVDLA_CSC_dl_for_check.scala 646:47:@811.4]
  assign _T_1072 = _GEN_712 * h_bias_3_stride; // @[NV_NVDLA_CSC_dl_for_check.scala 646:47:@811.4]
  assign _T_1073 = layer_st ? 19'h0 : _T_1072; // @[NV_NVDLA_CSC_dl_for_check.scala 646:21:@812.4]
  assign h_bias_3_w = _T_1073[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 646:65:@813.4]
  assign _T_1074 = is_winograd_d1[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 647:69:@814.4]
  assign _T_1075 = is_img_d1[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 647:84:@815.4]
  assign _T_1076 = _T_1074 | _T_1075; // @[NV_NVDLA_CSC_dl_for_check.scala 647:73:@816.4]
  assign _T_1077 = dat_exec_valid & _T_1076; // @[NV_NVDLA_CSC_dl_for_check.scala 647:52:@817.4]
  assign _T_1078 = layer_st | _T_1077; // @[NV_NVDLA_CSC_dl_for_check.scala 647:34:@818.4]
  assign h_bias_reg_en = {_T_1078,dat_exec_valid}; // @[Cat.scala 30:58:@819.4]
  assign _GEN_93 = datain_c_cnt_reg_en ? c_bias_w : c_bias; // @[NV_NVDLA_CSC_dl_for_check.scala 677:20:@840.4]
  assign _GEN_94 = c_bias_d1_reg_en ? c_bias : c_bias_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 680:23:@843.4]
  assign _T_1101 = h_bias_reg_en[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 683:19:@846.4]
  assign _GEN_95 = _T_1101 ? h_bias_0_w : h_bias_0_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 683:23:@847.4]
  assign _GEN_96 = _T_1101 ? h_bias_1_w : h_bias_1_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 683:23:@847.4]
  assign _GEN_97 = _T_1101 ? h_bias_2_w : h_bias_2_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 683:23:@847.4]
  assign _T_1102 = h_bias_reg_en[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 688:19:@852.4]
  assign _GEN_98 = _T_1102 ? h_bias_3_w : h_bias_3_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 688:23:@853.4]
  assign _GEN_99 = dat_exec_valid ? w_bias_w : {{1'd0}, w_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 691:20:@856.4]
  assign _T_1197 = h_bias_0_d1 + h_bias_1_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 717:30:@886.4]
  assign _GEN_713 = {{1'd0}, h_bias_2_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 717:45:@887.4]
  assign _T_1198 = _T_1197 + _GEN_713; // @[NV_NVDLA_CSC_dl_for_check.scala 717:45:@887.4]
  assign _GEN_714 = {{2'd0}, h_bias_3_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 717:60:@888.4]
  assign _T_1199 = _T_1198 + _GEN_714; // @[NV_NVDLA_CSC_dl_for_check.scala 717:60:@888.4]
  assign h_bias_d1 = _T_1199[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 717:75:@889.4]
  assign _GEN_715 = {{2'd0}, c_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 718:40:@890.4]
  assign _T_1200 = dat_entry_st + _GEN_715; // @[NV_NVDLA_CSC_dl_for_check.scala 718:40:@890.4]
  assign _GEN_716 = {{3'd0}, h_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 718:53:@891.4]
  assign _T_1201 = _T_1200 + _GEN_716; // @[NV_NVDLA_CSC_dl_for_check.scala 718:53:@891.4]
  assign _GEN_717 = {{4'd0}, w_bias_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 718:66:@892.4]
  assign dat_req_addr_sum = _T_1201 + _GEN_717; // @[NV_NVDLA_CSC_dl_for_check.scala 718:66:@892.4]
  assign _GEN_718 = {{3'd0}, _T_606}; // @[NV_NVDLA_CSC_dl_for_check.scala 719:45:@895.4]
  assign is_dat_req_addr_wrap = dat_req_addr_sum >= _GEN_718; // @[NV_NVDLA_CSC_dl_for_check.scala 719:45:@895.4]
  assign _T_1214 = dat_req_addr_sum - _GEN_718; // @[NV_NVDLA_CSC_dl_for_check.scala 720:42:@898.4]
  assign dat_req_addr_wrap = $unsigned(_T_1214); // @[NV_NVDLA_CSC_dl_for_check.scala 720:42:@899.4]
  assign _T_1215 = layer_st | dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 721:35:@900.4]
  assign _T_1221 = is_dat_req_addr_wrap ? dat_req_addr_wrap : {{1'd0}, dat_req_addr_sum}; // @[NV_NVDLA_CSC_dl_for_check.scala 722:25:@902.4]
  assign dat_req_addr_w = _T_1215 ? 19'h1fff : _T_1221; // @[NV_NVDLA_CSC_dl_for_check.scala 721:25:@903.4]
  assign _T_1225 = 2'h2 == dat_req_sub_h_d1; // @[Mux.scala 46:19:@904.4]
  assign _T_1226 = _T_1225 ? dat_req_sub_h_addr_2 : dat_req_sub_h_addr_3; // @[Mux.scala 46:16:@905.4]
  assign _T_1227 = 2'h1 == dat_req_sub_h_d1; // @[Mux.scala 46:19:@906.4]
  assign _T_1228 = _T_1227 ? dat_req_sub_h_addr_1 : _T_1226; // @[Mux.scala 46:16:@907.4]
  assign _T_1229 = 2'h0 == dat_req_sub_h_d1; // @[Mux.scala 46:19:@908.4]
  assign dat_req_addr_last = _T_1229 ? dat_req_sub_h_addr_0 : _T_1228; // @[Mux.scala 46:16:@909.4]
  assign _GEN_720 = {{6'd0}, dat_req_addr_last}; // @[NV_NVDLA_CSC_dl_for_check.scala 725:65:@910.4]
  assign _T_1230 = _GEN_720 != dat_req_addr_w; // @[NV_NVDLA_CSC_dl_for_check.scala 725:65:@910.4]
  assign _T_1231 = _T_1230 | pixel_force_fetch_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 725:85:@911.4]
  assign sc2buf_dat_rd_en_w = dat_req_valid_d1 & _T_1231; // @[NV_NVDLA_CSC_dl_for_check.scala 725:43:@912.4]
  assign _T_1232 = dat_req_valid_d1 | dat_req_dummy_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 727:38:@913.4]
  assign _T_1234 = dat_req_sub_h_d1 == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@914.4]
  assign _T_1235 = _T_1232 & _T_1234; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@915.4]
  assign dat_req_sub_h_addr_en_0 = layer_st | _T_1235; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@916.4]
  assign _T_1239 = dat_req_sub_h_d1 == 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@918.4]
  assign _T_1240 = _T_1232 & _T_1239; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@919.4]
  assign dat_req_sub_h_addr_en_1 = layer_st | _T_1240; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@920.4]
  assign _T_1244 = dat_req_sub_h_d1 == 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@922.4]
  assign _T_1245 = _T_1232 & _T_1244; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@923.4]
  assign dat_req_sub_h_addr_en_2 = layer_st | _T_1245; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@924.4]
  assign _T_1249 = dat_req_sub_h_d1 == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 727:78:@926.4]
  assign _T_1250 = _T_1232 & _T_1249; // @[NV_NVDLA_CSC_dl_for_check.scala 727:58:@927.4]
  assign dat_req_sub_h_addr_en_3 = layer_st | _T_1250; // @[NV_NVDLA_CSC_dl_for_check.scala 727:17:@928.4]
  assign _GEN_100 = dat_req_sub_h_addr_en_0 ? dat_req_addr_w : {{6'd0}, dat_req_sub_h_addr_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@934.4]
  assign _GEN_101 = dat_req_sub_h_addr_en_1 ? dat_req_addr_w : {{6'd0}, dat_req_sub_h_addr_1}; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@937.4]
  assign _GEN_102 = dat_req_sub_h_addr_en_2 ? dat_req_addr_w : {{6'd0}, dat_req_sub_h_addr_2}; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@940.4]
  assign _GEN_103 = dat_req_sub_h_addr_en_3 ? dat_req_addr_w : {{6'd0}, dat_req_sub_h_addr_3}; // @[NV_NVDLA_CSC_dl_for_check.scala 734:35:@943.4]
  assign _T_1261 = layer_st | sc2buf_dat_rd_en_w; // @[NV_NVDLA_CSC_dl_for_check.scala 740:14:@947.4]
  assign _GEN_104 = _T_1261 ? dat_req_addr_w : sc2buf_dat_rd_addr_out; // @[NV_NVDLA_CSC_dl_for_check.scala 740:34:@948.4]
  assign _GEN_105 = dat_exec_valid_d1 ? dat_req_sub_w_d1 : dat_req_pipe_sub_w; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_106 = dat_exec_valid_d1 ? dat_req_sub_h_d1 : dat_req_pipe_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_107 = dat_exec_valid_d1 ? dat_req_sub_c_d1 : dat_req_pipe_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_108 = dat_exec_valid_d1 ? dat_req_ch_end_d1 : dat_req_pipe_ch_end; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_109 = dat_exec_valid_d1 ? dat_req_bytes_d1 : dat_req_pipe_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_110 = dat_exec_valid_d1 ? dat_req_dummy_d1 : dat_req_pipe_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_111 = dat_exec_valid_d1 ? dat_req_cur_sub_h_d1 : dat_req_pipe_cur_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_112 = dat_exec_valid_d1 ? dat_req_sub_w_st_d1 : dat_req_pipe_sub_w_st; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_113 = dat_exec_valid_d1 ? dat_req_rls_d1 : dat_req_pipe_rls; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_114 = dat_exec_valid_d1 ? dat_req_flag_d1 : dat_req_pipe_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _GEN_115 = dat_exec_valid_d1 ? dat_req_dummy_d1 : dat_req_exec_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 748:24:@955.4]
  assign _T_1266 = {1'h0,dat_req_pipe_ch_end,dat_req_pipe_sub_c,dat_req_pipe_sub_h,dat_req_pipe_sub_w}; // @[Cat.scala 30:58:@971.4]
  assign dat_req_pipe_pd = {dat_req_pipe_flag,dat_req_pipe_rls,dat_req_pipe_sub_w_st,dat_req_pipe_dummy,dat_req_pipe_cur_sub_h,dat_req_pipe_bytes,_T_1266}; // @[Cat.scala 30:58:@977.4]
  assign _GEN_116 = dat_req_pipe_pvld ? dat_req_pipe_pd : _T_1295; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1019.4]
  assign _GEN_117 = dat_req_exec_pvld ? dat_req_exec_dummy : _T_1333; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1023.4]
  assign _GEN_118 = dat_req_exec_pvld ? 2'h0 : _T_1352; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1023.4]
  assign _GEN_119 = _T_1276 ? _T_1295 : _T_1298; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1028.4]
  assign _GEN_120 = _T_1314 ? _T_1333 : _T_1336; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1032.4]
  assign _GEN_121 = _T_1314 ? _T_1352 : _T_1355; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1032.4]
  assign _GEN_122 = _T_1279 ? _T_1298 : _T_1301; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1037.4]
  assign _GEN_123 = _T_1317 ? _T_1336 : _T_1339; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1041.4]
  assign _GEN_124 = _T_1317 ? _T_1355 : _T_1358; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1041.4]
  assign _GEN_125 = _T_1282 ? _T_1301 : _T_1304; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1046.4]
  assign _GEN_126 = _T_1320 ? _T_1339 : _T_1342; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1050.4]
  assign _GEN_127 = _T_1320 ? _T_1358 : _T_1361; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1050.4]
  assign _GEN_128 = _T_1285 ? _T_1304 : _T_1307; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1055.4]
  assign _GEN_129 = _T_1323 ? _T_1342 : _T_1345; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1059.4]
  assign _GEN_130 = _T_1323 ? _T_1361 : _T_1364; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1059.4]
  assign _GEN_131 = _T_1288 ? _T_1307 : dat_rsp_pipe_pd; // @[NV_NVDLA_CSC_dl_for_check.scala 792:33:@1064.4]
  assign _GEN_132 = _T_1326 ? _T_1345 : dat_rsp_exec_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1068.4]
  assign _GEN_133 = _T_1326 ? _T_1364 : dat_rsp_exec_sub_h; // @[NV_NVDLA_CSC_dl_for_check.scala 796:33:@1068.4]
  assign dat_rsp_pipe_sub_w = dat_rsp_pipe_pd[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 809:41:@1072.4]
  assign dat_rsp_pipe_sub_h = dat_rsp_pipe_pd[3:2]; // @[NV_NVDLA_CSC_dl_for_check.scala 810:41:@1073.4]
  assign dat_rsp_pipe_sub_c = dat_rsp_pipe_pd[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 811:41:@1074.4]
  assign dat_rsp_pipe_ch_end = dat_rsp_pipe_pd[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 812:42:@1075.4]
  assign dat_rsp_pipe_bytes = dat_rsp_pipe_pd[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 813:41:@1076.4]
  assign dat_rsp_pipe_cur_sub_h = dat_rsp_pipe_pd[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 814:45:@1077.4]
  assign dat_rsp_pipe_sub_w_st = dat_rsp_pipe_pd[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 816:44:@1079.4]
  assign dat_rsp_pipe_rls = dat_rsp_pipe_pd[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 817:39:@1080.4]
  assign dat_rsp_pipe_flag = dat_rsp_pipe_pd[28:20]; // @[NV_NVDLA_CSC_dl_for_check.scala 818:40:@1081.4]
  assign _T_1392 = dat_rsp_exec_sub_h == 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 841:70:@1098.4]
  assign dat_l0c0_en = io_sc2buf_dat_rd_data_valid & _T_1392; // @[NV_NVDLA_CSC_dl_for_check.scala 841:48:@1099.4]
  assign _T_1394 = dat_rsp_exec_sub_h == 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 842:70:@1100.4]
  assign dat_l1c0_en = io_sc2buf_dat_rd_data_valid & _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 842:48:@1101.4]
  assign _T_1396 = dat_rsp_exec_sub_h == 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 843:70:@1102.4]
  assign dat_l2c0_en = io_sc2buf_dat_rd_data_valid & _T_1396; // @[NV_NVDLA_CSC_dl_for_check.scala 843:48:@1103.4]
  assign _T_1398 = dat_rsp_exec_sub_h == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 844:70:@1104.4]
  assign dat_l3c0_en = io_sc2buf_dat_rd_data_valid & _T_1398; // @[NV_NVDLA_CSC_dl_for_check.scala 844:48:@1105.4]
  assign _T_1399 = is_winograd_d1[11]; // @[NV_NVDLA_CSC_dl_for_check.scala 847:62:@1106.4]
  assign _T_1400 = io_sc2buf_dat_rd_data_valid & _T_1399; // @[NV_NVDLA_CSC_dl_for_check.scala 847:46:@1107.4]
  assign _T_1401 = ~ dat_rsp_pipe_sub_w_st; // @[NV_NVDLA_CSC_dl_for_check.scala 847:69:@1108.4]
  assign dat_wg_adv = _T_1400 & _T_1401; // @[NV_NVDLA_CSC_dl_for_check.scala 847:67:@1109.4]
  assign _T_1402 = dat_rsp_exec_sub_h[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 848:52:@1110.4]
  assign _T_1403 = ~ _T_1402; // @[NV_NVDLA_CSC_dl_for_check.scala 848:33:@1111.4]
  assign _T_1404 = dat_wg_adv & _T_1403; // @[NV_NVDLA_CSC_dl_for_check.scala 848:31:@1112.4]
  assign _T_1405 = is_img_d1[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 848:69:@1113.4]
  assign _T_1406 = _T_1405 & dat_l0c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 848:74:@1114.4]
  assign _T_1407 = ~ dat_l0c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 848:90:@1115.4]
  assign _T_1408 = _T_1406 & _T_1407; // @[NV_NVDLA_CSC_dl_for_check.scala 848:88:@1116.4]
  assign dat_l0c1_en = _T_1404 | _T_1408; // @[NV_NVDLA_CSC_dl_for_check.scala 848:57:@1117.4]
  assign _T_1410 = dat_wg_adv & _T_1402; // @[NV_NVDLA_CSC_dl_for_check.scala 849:31:@1119.4]
  assign _T_1411 = is_img_d1[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 849:68:@1120.4]
  assign _T_1412 = _T_1411 & dat_l1c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 849:73:@1121.4]
  assign _T_1413 = ~ dat_l1c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 849:89:@1122.4]
  assign _T_1414 = _T_1412 & _T_1413; // @[NV_NVDLA_CSC_dl_for_check.scala 849:87:@1123.4]
  assign dat_l1c1_en = _T_1410 | _T_1414; // @[NV_NVDLA_CSC_dl_for_check.scala 849:56:@1124.4]
  assign _T_1415 = is_img_d1[15]; // @[NV_NVDLA_CSC_dl_for_check.scala 850:29:@1125.4]
  assign _T_1416 = _T_1415 & dat_l2c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 850:34:@1126.4]
  assign _T_1417 = ~ dat_l2c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 850:50:@1127.4]
  assign dat_l2c1_en = _T_1416 & _T_1417; // @[NV_NVDLA_CSC_dl_for_check.scala 850:48:@1128.4]
  assign _T_1418 = is_img_d1[16]; // @[NV_NVDLA_CSC_dl_for_check.scala 851:29:@1129.4]
  assign _T_1419 = _T_1418 & dat_l3c0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 851:34:@1130.4]
  assign _T_1420 = ~ dat_l3c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 851:50:@1131.4]
  assign dat_l3c1_en = _T_1419 & _T_1420; // @[NV_NVDLA_CSC_dl_for_check.scala 851:48:@1132.4]
  assign _T_1421 = dat_rsp_exec_pvld & dat_rsp_exec_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 853:41:@1133.4]
  assign dat_dummy_l0_en = _T_1421 & _T_1392; // @[NV_NVDLA_CSC_dl_for_check.scala 853:62:@1135.4]
  assign dat_dummy_l1_en = _T_1421 & _T_1394; // @[NV_NVDLA_CSC_dl_for_check.scala 854:62:@1138.4]
  assign dat_dummy_l2_en = _T_1421 & _T_1396; // @[NV_NVDLA_CSC_dl_for_check.scala 855:62:@1141.4]
  assign dat_dummy_l3_en = _T_1421 & _T_1398; // @[NV_NVDLA_CSC_dl_for_check.scala 856:62:@1144.4]
  assign dat_l0_set = dat_l0c0_en | dat_dummy_l0_en; // @[NV_NVDLA_CSC_dl_for_check.scala 858:30:@1145.4]
  assign dat_l1_set = dat_l1c0_en | dat_dummy_l1_en; // @[NV_NVDLA_CSC_dl_for_check.scala 859:30:@1146.4]
  assign dat_l2_set = dat_l2c0_en | dat_dummy_l2_en; // @[NV_NVDLA_CSC_dl_for_check.scala 860:30:@1147.4]
  assign dat_l3_set = dat_l3c0_en | dat_dummy_l3_en; // @[NV_NVDLA_CSC_dl_for_check.scala 861:30:@1148.4]
  assign _T_1435 = dat_dummy_l0_en ? 1'h1 : dat_l0c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 863:48:@1149.4]
  assign _T_1436 = dat_l0c0_en ? 1'h0 : _T_1435; // @[NV_NVDLA_CSC_dl_for_check.scala 863:22:@1150.4]
  assign _T_1439 = dat_dummy_l1_en ? 1'h1 : dat_l1c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 864:48:@1152.4]
  assign _T_1440 = dat_l1c0_en ? 1'h0 : _T_1439; // @[NV_NVDLA_CSC_dl_for_check.scala 864:22:@1153.4]
  assign _T_1443 = dat_dummy_l2_en ? 1'h1 : dat_l2c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 865:48:@1155.4]
  assign _T_1444 = dat_l2c0_en ? 1'h0 : _T_1443; // @[NV_NVDLA_CSC_dl_for_check.scala 865:22:@1156.4]
  assign _T_1447 = dat_dummy_l3_en ? 1'h1 : dat_l3c0_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 866:48:@1158.4]
  assign _T_1448 = dat_l3c0_en ? 1'h0 : _T_1447; // @[NV_NVDLA_CSC_dl_for_check.scala 866:22:@1159.4]
  assign _T_1450 = dat_l0_set ? dat_l0c0_dummy : dat_l0c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 867:48:@1161.4]
  assign _T_1451 = dat_l0c1_en ? 1'h0 : _T_1450; // @[NV_NVDLA_CSC_dl_for_check.scala 867:22:@1162.4]
  assign _T_1454 = sub_h_total_g2 != 2'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 868:77:@1164.4]
  assign _T_1455 = dat_l1_set & _T_1454; // @[NV_NVDLA_CSC_dl_for_check.scala 868:60:@1165.4]
  assign _T_1456 = _T_1455 ? dat_l1c0_dummy : dat_l1c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 868:48:@1166.4]
  assign _T_1457 = dat_l1c1_en ? 1'h0 : _T_1456; // @[NV_NVDLA_CSC_dl_for_check.scala 868:22:@1167.4]
  assign _T_1459 = sub_h_total_g2[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 869:76:@1169.4]
  assign _T_1460 = dat_l2_set & _T_1459; // @[NV_NVDLA_CSC_dl_for_check.scala 869:60:@1170.4]
  assign _T_1461 = _T_1460 ? dat_l2c0_dummy : dat_l2c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 869:48:@1171.4]
  assign _T_1462 = dat_l2c1_en ? 1'h0 : _T_1461; // @[NV_NVDLA_CSC_dl_for_check.scala 869:22:@1172.4]
  assign _T_1465 = dat_l3_set & _T_1459; // @[NV_NVDLA_CSC_dl_for_check.scala 870:60:@1175.4]
  assign _T_1466 = _T_1465 ? dat_l3c0_dummy : dat_l3c1_dummy; // @[NV_NVDLA_CSC_dl_for_check.scala 870:48:@1176.4]
  assign _T_1467 = dat_l3c1_en ? 1'h0 : _T_1466; // @[NV_NVDLA_CSC_dl_for_check.scala 870:22:@1177.4]
  assign _T_1516 = {dat_rsp_pipe_flag,dat_rsp_pipe_rls,dat_rsp_pipe_cur_sub_h,dat_rsp_pipe_bytes,1'h0,dat_rsp_pipe_ch_end,dat_rsp_pipe_sub_c,dat_rsp_pipe_sub_h,dat_rsp_pipe_sub_w}; // @[Cat.scala 30:58:@1229.4]
  assign _GEN_142 = dat_rsp_pipe_pvld ? _T_1516 : _T_1498; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1232.4]
  assign _GEN_143 = dat_rsp_l0_pvld ? _T_1498 : _T_1501; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1236.4]
  assign _GEN_144 = dat_rsp_l1_pvld ? _T_1501 : _T_1504; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1240.4]
  assign _GEN_145 = dat_rsp_l2_pvld ? _T_1504 : _T_1507; // @[NV_NVDLA_CSC_dl_for_check.scala 906:28:@1244.4]
  assign dat_rsp_l0_sub_c = _T_1498[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 924:39:@1270.4]
  assign dat_rsp_l1_sub_c = _T_1501[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 925:39:@1271.4]
  assign dat_rsp_l2_sub_c = _T_1504[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 926:39:@1272.4]
  assign dat_rsp_l3_sub_c = _T_1507[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 927:39:@1273.4]
  assign dat_rsp_l0_flag = _T_1498[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 929:38:@1274.4]
  assign dat_rsp_l1_flag = _T_1501[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 930:38:@1275.4]
  assign dat_rsp_l2_flag = _T_1504[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 931:38:@1276.4]
  assign dat_rsp_l3_flag = _T_1507[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 932:38:@1277.4]
  assign dat_rsp_l0_stripe_end = dat_rsp_l0_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 934:44:@1278.4]
  assign dat_rsp_l1_stripe_end = dat_rsp_l1_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 935:44:@1279.4]
  assign dat_rsp_l2_stripe_end = dat_rsp_l2_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 936:44:@1280.4]
  assign dat_rsp_l3_stripe_end = dat_rsp_l3_flag[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 937:44:@1281.4]
  assign dat_rsp_sub_w = dat_rsp_pd[1:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 940:31:@1282.4]
  assign dat_rsp_bytes = dat_rsp_pd[14:7]; // @[NV_NVDLA_CSC_dl_for_check.scala 944:31:@1286.4]
  assign dat_rsp_cur_sub_h = dat_rsp_pd[16:15]; // @[NV_NVDLA_CSC_dl_for_check.scala 945:35:@1287.4]
  assign dat_rsp_flag = dat_rsp_pd[26:18]; // @[NV_NVDLA_CSC_dl_for_check.scala 947:30:@1290.4]
  assign rsp_sft_cnt_l0_sub = dat_l0c0_en ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 956:29:@1296.4]
  assign rsp_sft_cnt_l1_sub = dat_l1c0_en ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 957:29:@1297.4]
  assign rsp_sft_cnt_l2_sub = dat_l2c0_en ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 958:29:@1298.4]
  assign rsp_sft_cnt_l3_sub = dat_l3c0_en ? 8'h40 : 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 959:29:@1299.4]
  assign _T_1554 = pixel_x_byte_stride > 7'h40; // @[NV_NVDLA_CSC_dl_for_check.scala 961:50:@1300.4]
  assign _GEN_721 = {{1'd0}, pixel_x_byte_stride}; // @[NV_NVDLA_CSC_dl_for_check.scala 961:111:@1301.4]
  assign _T_1556 = rsp_sft_cnt_l0 + _GEN_721; // @[NV_NVDLA_CSC_dl_for_check.scala 961:111:@1301.4]
  assign _GEN_722 = {{1'd0}, rsp_sft_cnt_l0_sub}; // @[NV_NVDLA_CSC_dl_for_check.scala 961:134:@1302.4]
  assign _T_1557 = _T_1556 - _GEN_722; // @[NV_NVDLA_CSC_dl_for_check.scala 961:134:@1302.4]
  assign _T_1558 = $unsigned(_T_1557); // @[NV_NVDLA_CSC_dl_for_check.scala 961:134:@1303.4]
  assign _T_1559 = _T_1554 ? 10'h40 : _T_1558; // @[NV_NVDLA_CSC_dl_for_check.scala 961:29:@1304.4]
  assign rsp_sft_cnt_l0_inc = _T_1559[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 961:156:@1305.4]
  assign _T_1563 = rsp_sft_cnt_l1 + _GEN_721; // @[NV_NVDLA_CSC_dl_for_check.scala 962:111:@1307.4]
  assign _GEN_724 = {{1'd0}, rsp_sft_cnt_l1_sub}; // @[NV_NVDLA_CSC_dl_for_check.scala 962:134:@1308.4]
  assign _T_1564 = _T_1563 - _GEN_724; // @[NV_NVDLA_CSC_dl_for_check.scala 962:134:@1308.4]
  assign _T_1565 = $unsigned(_T_1564); // @[NV_NVDLA_CSC_dl_for_check.scala 962:134:@1309.4]
  assign _T_1566 = _T_1554 ? 10'h40 : _T_1565; // @[NV_NVDLA_CSC_dl_for_check.scala 962:29:@1310.4]
  assign rsp_sft_cnt_l1_inc = _T_1566[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 962:156:@1311.4]
  assign _T_1570 = rsp_sft_cnt_l2 + _GEN_721; // @[NV_NVDLA_CSC_dl_for_check.scala 963:111:@1313.4]
  assign _GEN_726 = {{1'd0}, rsp_sft_cnt_l2_sub}; // @[NV_NVDLA_CSC_dl_for_check.scala 963:134:@1314.4]
  assign _T_1571 = _T_1570 - _GEN_726; // @[NV_NVDLA_CSC_dl_for_check.scala 963:134:@1314.4]
  assign _T_1572 = $unsigned(_T_1571); // @[NV_NVDLA_CSC_dl_for_check.scala 963:134:@1315.4]
  assign _T_1573 = _T_1554 ? 10'h40 : _T_1572; // @[NV_NVDLA_CSC_dl_for_check.scala 963:29:@1316.4]
  assign rsp_sft_cnt_l2_inc = _T_1573[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 963:156:@1317.4]
  assign _T_1577 = rsp_sft_cnt_l3 + _GEN_721; // @[NV_NVDLA_CSC_dl_for_check.scala 964:111:@1319.4]
  assign _GEN_728 = {{1'd0}, rsp_sft_cnt_l3_sub}; // @[NV_NVDLA_CSC_dl_for_check.scala 964:134:@1320.4]
  assign _T_1578 = _T_1577 - _GEN_728; // @[NV_NVDLA_CSC_dl_for_check.scala 964:134:@1320.4]
  assign _T_1579 = $unsigned(_T_1578); // @[NV_NVDLA_CSC_dl_for_check.scala 964:134:@1321.4]
  assign _T_1580 = _T_1554 ? 10'h40 : _T_1579; // @[NV_NVDLA_CSC_dl_for_check.scala 964:29:@1322.4]
  assign rsp_sft_cnt_l3_inc = _T_1580[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 964:156:@1323.4]
  assign _T_1582 = ~ dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 973:52:@1324.4]
  assign _T_1583 = dat_rsp_l0_stripe_end & _T_1582; // @[NV_NVDLA_CSC_dl_for_check.scala 973:50:@1325.4]
  assign _T_1584 = dat_rsp_l0_stripe_end & dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 974:50:@1326.4]
  assign _T_1587 = rsp_sft_cnt_l0_inc & 8'h3f; // @[NV_NVDLA_CSC_dl_for_check.scala 975:64:@1327.4]
  assign _T_1588 = dat_dummy_l0_en ? _T_1587 : rsp_sft_cnt_l0_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 975:27:@1328.4]
  assign _T_1589 = _T_1584 ? 8'h40 : _T_1588; // @[NV_NVDLA_CSC_dl_for_check.scala 974:27:@1329.4]
  assign _T_1590 = _T_1583 ? rsp_sft_cnt_l0_ori : _T_1589; // @[NV_NVDLA_CSC_dl_for_check.scala 973:27:@1330.4]
  assign rsp_sft_cnt_l0_w = layer_st ? 8'h40 : _T_1590; // @[NV_NVDLA_CSC_dl_for_check.scala 972:27:@1331.4]
  assign _T_1592 = ~ dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 978:52:@1332.4]
  assign _T_1593 = dat_rsp_l1_stripe_end & _T_1592; // @[NV_NVDLA_CSC_dl_for_check.scala 978:50:@1333.4]
  assign _T_1594 = dat_rsp_l1_stripe_end & dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 979:50:@1334.4]
  assign _T_1597 = rsp_sft_cnt_l1_inc & 8'h3f; // @[NV_NVDLA_CSC_dl_for_check.scala 980:64:@1335.4]
  assign _T_1598 = dat_dummy_l1_en ? _T_1597 : rsp_sft_cnt_l1_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 980:27:@1336.4]
  assign _T_1599 = _T_1594 ? 8'h40 : _T_1598; // @[NV_NVDLA_CSC_dl_for_check.scala 979:27:@1337.4]
  assign _T_1600 = _T_1593 ? rsp_sft_cnt_l1_ori : _T_1599; // @[NV_NVDLA_CSC_dl_for_check.scala 978:27:@1338.4]
  assign rsp_sft_cnt_l1_w = layer_st ? 8'h40 : _T_1600; // @[NV_NVDLA_CSC_dl_for_check.scala 977:27:@1339.4]
  assign _T_1602 = ~ dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 983:52:@1340.4]
  assign _T_1603 = dat_rsp_l2_stripe_end & _T_1602; // @[NV_NVDLA_CSC_dl_for_check.scala 983:50:@1341.4]
  assign _T_1604 = dat_rsp_l2_stripe_end & dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 984:50:@1342.4]
  assign _T_1607 = rsp_sft_cnt_l2_inc & 8'h3f; // @[NV_NVDLA_CSC_dl_for_check.scala 985:64:@1343.4]
  assign _T_1608 = dat_dummy_l2_en ? _T_1607 : rsp_sft_cnt_l2_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 985:27:@1344.4]
  assign _T_1609 = _T_1604 ? 8'h40 : _T_1608; // @[NV_NVDLA_CSC_dl_for_check.scala 984:27:@1345.4]
  assign _T_1610 = _T_1603 ? rsp_sft_cnt_l2_ori : _T_1609; // @[NV_NVDLA_CSC_dl_for_check.scala 983:27:@1346.4]
  assign rsp_sft_cnt_l2_w = layer_st ? 8'h40 : _T_1610; // @[NV_NVDLA_CSC_dl_for_check.scala 982:27:@1347.4]
  assign _T_1612 = ~ dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 988:52:@1348.4]
  assign _T_1613 = dat_rsp_l3_stripe_end & _T_1612; // @[NV_NVDLA_CSC_dl_for_check.scala 988:50:@1349.4]
  assign _T_1614 = dat_rsp_l3_stripe_end & dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 989:50:@1350.4]
  assign _T_1617 = rsp_sft_cnt_l3_inc & 8'h3f; // @[NV_NVDLA_CSC_dl_for_check.scala 990:64:@1351.4]
  assign _T_1618 = dat_dummy_l3_en ? _T_1617 : rsp_sft_cnt_l3_inc; // @[NV_NVDLA_CSC_dl_for_check.scala 990:27:@1352.4]
  assign _T_1619 = _T_1614 ? 8'h40 : _T_1618; // @[NV_NVDLA_CSC_dl_for_check.scala 989:27:@1353.4]
  assign _T_1620 = _T_1613 ? rsp_sft_cnt_l3_ori : _T_1619; // @[NV_NVDLA_CSC_dl_for_check.scala 988:27:@1354.4]
  assign rsp_sft_cnt_l3_w = layer_st ? 8'h40 : _T_1620; // @[NV_NVDLA_CSC_dl_for_check.scala 987:27:@1355.4]
  assign _T_1621 = is_img_d1[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 993:46:@1356.4]
  assign _T_1622 = _T_1621 & dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 993:51:@1357.4]
  assign rsp_sft_cnt_l0_en = layer_st | _T_1622; // @[NV_NVDLA_CSC_dl_for_check.scala 993:34:@1358.4]
  assign _T_1623 = is_img_d1[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 994:46:@1359.4]
  assign _T_1624 = _T_1623 & dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 994:51:@1360.4]
  assign _T_1626 = sub_h_total_g5 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 994:87:@1361.4]
  assign _T_1627 = _T_1624 & _T_1626; // @[NV_NVDLA_CSC_dl_for_check.scala 994:69:@1362.4]
  assign rsp_sft_cnt_l1_en = layer_st | _T_1627; // @[NV_NVDLA_CSC_dl_for_check.scala 994:34:@1363.4]
  assign _T_1628 = is_img_d1[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 995:46:@1364.4]
  assign _T_1629 = _T_1628 & dat_rsp_l2_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 995:51:@1365.4]
  assign _T_1631 = sub_h_total_g5 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 995:87:@1366.4]
  assign _T_1632 = _T_1629 & _T_1631; // @[NV_NVDLA_CSC_dl_for_check.scala 995:69:@1367.4]
  assign rsp_sft_cnt_l2_en = layer_st | _T_1632; // @[NV_NVDLA_CSC_dl_for_check.scala 995:34:@1368.4]
  assign _T_1633 = is_img_d1[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 996:46:@1369.4]
  assign _T_1634 = _T_1633 & dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 996:51:@1370.4]
  assign _T_1637 = _T_1634 & _T_1631; // @[NV_NVDLA_CSC_dl_for_check.scala 996:69:@1372.4]
  assign rsp_sft_cnt_l3_en = layer_st | _T_1637; // @[NV_NVDLA_CSC_dl_for_check.scala 996:34:@1373.4]
  assign _T_1638 = is_img_d1[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 998:50:@1374.4]
  assign _T_1639 = _T_1638 & dat_rsp_l0_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 998:55:@1375.4]
  assign _T_1640 = _T_1639 & dat_rsp_l0_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 998:73:@1376.4]
  assign _T_1641 = _T_1640 & dat_rsp_l0_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 998:97:@1377.4]
  assign rsp_sft_cnt_l0_ori_en = layer_st | _T_1641; // @[NV_NVDLA_CSC_dl_for_check.scala 998:38:@1378.4]
  assign _T_1642 = is_img_d1[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 999:50:@1379.4]
  assign _T_1643 = _T_1642 & dat_rsp_l1_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 999:55:@1380.4]
  assign _T_1644 = _T_1643 & dat_rsp_l1_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 999:73:@1381.4]
  assign _T_1645 = _T_1644 & dat_rsp_l1_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 999:97:@1382.4]
  assign _T_1647 = sub_h_total_g6 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 999:138:@1383.4]
  assign _T_1648 = _T_1645 & _T_1647; // @[NV_NVDLA_CSC_dl_for_check.scala 999:120:@1384.4]
  assign rsp_sft_cnt_l1_ori_en = layer_st | _T_1648; // @[NV_NVDLA_CSC_dl_for_check.scala 999:38:@1385.4]
  assign _T_1649 = is_img_d1[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:50:@1386.4]
  assign _T_1650 = _T_1649 & dat_rsp_l2_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:55:@1387.4]
  assign _T_1651 = _T_1650 & dat_rsp_l2_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:73:@1388.4]
  assign _T_1652 = _T_1651 & dat_rsp_l2_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:97:@1389.4]
  assign _T_1654 = sub_h_total_g6 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:138:@1390.4]
  assign _T_1655 = _T_1652 & _T_1654; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:120:@1391.4]
  assign rsp_sft_cnt_l2_ori_en = layer_st | _T_1655; // @[NV_NVDLA_CSC_dl_for_check.scala 1000:38:@1392.4]
  assign _T_1656 = is_img_d1[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:50:@1393.4]
  assign _T_1657 = _T_1656 & dat_rsp_l3_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:55:@1394.4]
  assign _T_1658 = _T_1657 & dat_rsp_l3_stripe_end; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:73:@1395.4]
  assign _T_1659 = _T_1658 & dat_rsp_l3_sub_c; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:97:@1396.4]
  assign _T_1662 = _T_1659 & _T_1654; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:120:@1398.4]
  assign rsp_sft_cnt_l3_ori_en = layer_st | _T_1662; // @[NV_NVDLA_CSC_dl_for_check.scala 1001:38:@1399.4]
  assign _GEN_146 = rsp_sft_cnt_l0_en ? rsp_sft_cnt_l0_w : rsp_sft_cnt_l0; // @[NV_NVDLA_CSC_dl_for_check.scala 1003:24:@1400.4]
  assign _GEN_147 = rsp_sft_cnt_l1_en ? rsp_sft_cnt_l1_w : rsp_sft_cnt_l1; // @[NV_NVDLA_CSC_dl_for_check.scala 1004:24:@1403.4]
  assign _GEN_148 = rsp_sft_cnt_l2_en ? rsp_sft_cnt_l2_w : rsp_sft_cnt_l2; // @[NV_NVDLA_CSC_dl_for_check.scala 1005:24:@1406.4]
  assign _GEN_149 = rsp_sft_cnt_l3_en ? rsp_sft_cnt_l3_w : rsp_sft_cnt_l3; // @[NV_NVDLA_CSC_dl_for_check.scala 1006:24:@1409.4]
  assign _GEN_150 = rsp_sft_cnt_l0_ori_en ? rsp_sft_cnt_l0_w : rsp_sft_cnt_l0_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1007:28:@1412.4]
  assign _GEN_151 = rsp_sft_cnt_l1_ori_en ? rsp_sft_cnt_l1_w : rsp_sft_cnt_l1_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1008:28:@1415.4]
  assign _GEN_152 = rsp_sft_cnt_l2_ori_en ? rsp_sft_cnt_l2_w : rsp_sft_cnt_l2_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1009:28:@1418.4]
  assign _GEN_153 = rsp_sft_cnt_l3_ori_en ? rsp_sft_cnt_l3_w : rsp_sft_cnt_l3_ori; // @[NV_NVDLA_CSC_dl_for_check.scala 1010:28:@1421.4]
  assign _T_1663 = pad_value[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1019:55:@1424.4]
  assign _T_1666 = {_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663}; // @[Cat.scala 30:58:@1427.4]
  assign _T_1667 = {_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1666}; // @[Cat.scala 30:58:@1428.4]
  assign _T_1668 = {_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1663,_T_1666,_T_1667}; // @[Cat.scala 30:58:@1429.4]
  assign dat_rsp_pad_value = {_T_1668,_T_1668}; // @[Cat.scala 30:58:@1430.4]
  assign dat_rsp_l0c0 = dat_l0c0_dummy ? dat_rsp_pad_value : dat_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1021:23:@1431.4]
  assign dat_rsp_l1c0 = dat_l1c0_dummy ? dat_rsp_pad_value : dat_l1c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1022:23:@1432.4]
  assign dat_rsp_l2c0 = dat_l2c0_dummy ? dat_rsp_pad_value : dat_l2c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1023:23:@1433.4]
  assign dat_rsp_l3c0 = dat_l3c0_dummy ? dat_rsp_pad_value : dat_l3c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1024:23:@1434.4]
  assign dat_rsp_l0c1 = dat_l0c1_dummy ? dat_rsp_pad_value : dat_l0c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1026:23:@1435.4]
  assign dat_rsp_l1c1 = dat_l1c1_dummy ? dat_rsp_pad_value : dat_l1c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1027:23:@1436.4]
  assign dat_rsp_l2c1 = dat_l2c1_dummy ? dat_rsp_pad_value : dat_l2c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1028:23:@1437.4]
  assign dat_rsp_l3c1 = dat_l3c1_dummy ? dat_rsp_pad_value : dat_l3c1; // @[NV_NVDLA_CSC_dl_for_check.scala 1029:23:@1438.4]
  assign _T_1670 = is_winograd_d1[14]; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:42:@1440.4]
  assign _T_1671 = is_img_d1[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:58:@1441.4]
  assign _T_1672 = _T_1670 | _T_1671; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:47:@1442.4]
  assign _T_1675 = dat_rsp_bytes <= 8'h20; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:43:@1443.4]
  assign _T_1676 = dat_rsp_sub_w[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:87:@1444.4]
  assign _T_1678 = _T_1676 == 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:91:@1445.4]
  assign _T_1679 = _T_1675 & _T_1678; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:72:@1446.4]
  assign _T_1681 = dat_rsp_l0c0[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:171:@1447.4]
  assign _T_1682 = {256'h0,_T_1681}; // @[Cat.scala 30:58:@1448.4]
  assign _T_1688 = _T_1675 & _T_1676; // @[NV_NVDLA_CSC_dl_for_check.scala 1041:72:@1452.4]
  assign _T_1690 = dat_rsp_l0c0[511:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1041:171:@1453.4]
  assign _T_1691 = {256'h0,_T_1690}; // @[Cat.scala 30:58:@1454.4]
  assign _T_1692 = _T_1688 ? _T_1691 : dat_rsp_l0c0; // @[NV_NVDLA_CSC_dl_for_check.scala 1041:27:@1455.4]
  assign _T_1693 = _T_1679 ? _T_1682 : _T_1692; // @[NV_NVDLA_CSC_dl_for_check.scala 1040:27:@1456.4]
  assign dat_rsp_conv_8b = _T_1672 ? 512'h0 : _T_1693; // @[NV_NVDLA_CSC_dl_for_check.scala 1039:27:@1457.4]
  assign dat_rsp_conv_0 = dat_rsp_conv_8b[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1460.4]
  assign dat_rsp_conv_1 = dat_rsp_conv_8b[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1462.4]
  assign dat_rsp_conv_2 = dat_rsp_conv_8b[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1464.4]
  assign dat_rsp_conv_3 = dat_rsp_conv_8b[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1466.4]
  assign dat_rsp_conv_4 = dat_rsp_conv_8b[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1468.4]
  assign dat_rsp_conv_5 = dat_rsp_conv_8b[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1470.4]
  assign dat_rsp_conv_6 = dat_rsp_conv_8b[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1472.4]
  assign dat_rsp_conv_7 = dat_rsp_conv_8b[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1474.4]
  assign dat_rsp_conv_8 = dat_rsp_conv_8b[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1476.4]
  assign dat_rsp_conv_9 = dat_rsp_conv_8b[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1478.4]
  assign dat_rsp_conv_10 = dat_rsp_conv_8b[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1480.4]
  assign dat_rsp_conv_11 = dat_rsp_conv_8b[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1482.4]
  assign dat_rsp_conv_12 = dat_rsp_conv_8b[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1484.4]
  assign dat_rsp_conv_13 = dat_rsp_conv_8b[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1486.4]
  assign dat_rsp_conv_14 = dat_rsp_conv_8b[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1488.4]
  assign dat_rsp_conv_15 = dat_rsp_conv_8b[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1490.4]
  assign dat_rsp_conv_16 = dat_rsp_conv_8b[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1492.4]
  assign dat_rsp_conv_17 = dat_rsp_conv_8b[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1494.4]
  assign dat_rsp_conv_18 = dat_rsp_conv_8b[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1496.4]
  assign dat_rsp_conv_19 = dat_rsp_conv_8b[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1498.4]
  assign dat_rsp_conv_20 = dat_rsp_conv_8b[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1500.4]
  assign dat_rsp_conv_21 = dat_rsp_conv_8b[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1502.4]
  assign dat_rsp_conv_22 = dat_rsp_conv_8b[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1504.4]
  assign dat_rsp_conv_23 = dat_rsp_conv_8b[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1506.4]
  assign dat_rsp_conv_24 = dat_rsp_conv_8b[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1508.4]
  assign dat_rsp_conv_25 = dat_rsp_conv_8b[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1510.4]
  assign dat_rsp_conv_26 = dat_rsp_conv_8b[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1512.4]
  assign dat_rsp_conv_27 = dat_rsp_conv_8b[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1514.4]
  assign dat_rsp_conv_28 = dat_rsp_conv_8b[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1516.4]
  assign dat_rsp_conv_29 = dat_rsp_conv_8b[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1518.4]
  assign dat_rsp_conv_30 = dat_rsp_conv_8b[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1520.4]
  assign dat_rsp_conv_31 = dat_rsp_conv_8b[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1522.4]
  assign dat_rsp_conv_32 = dat_rsp_conv_8b[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1524.4]
  assign dat_rsp_conv_33 = dat_rsp_conv_8b[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1526.4]
  assign dat_rsp_conv_34 = dat_rsp_conv_8b[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1528.4]
  assign dat_rsp_conv_35 = dat_rsp_conv_8b[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1530.4]
  assign dat_rsp_conv_36 = dat_rsp_conv_8b[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1532.4]
  assign dat_rsp_conv_37 = dat_rsp_conv_8b[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1534.4]
  assign dat_rsp_conv_38 = dat_rsp_conv_8b[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1536.4]
  assign dat_rsp_conv_39 = dat_rsp_conv_8b[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1538.4]
  assign dat_rsp_conv_40 = dat_rsp_conv_8b[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1540.4]
  assign dat_rsp_conv_41 = dat_rsp_conv_8b[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1542.4]
  assign dat_rsp_conv_42 = dat_rsp_conv_8b[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1544.4]
  assign dat_rsp_conv_43 = dat_rsp_conv_8b[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1546.4]
  assign dat_rsp_conv_44 = dat_rsp_conv_8b[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1548.4]
  assign dat_rsp_conv_45 = dat_rsp_conv_8b[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1550.4]
  assign dat_rsp_conv_46 = dat_rsp_conv_8b[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1552.4]
  assign dat_rsp_conv_47 = dat_rsp_conv_8b[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1554.4]
  assign dat_rsp_conv_48 = dat_rsp_conv_8b[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1556.4]
  assign dat_rsp_conv_49 = dat_rsp_conv_8b[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1558.4]
  assign dat_rsp_conv_50 = dat_rsp_conv_8b[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1560.4]
  assign dat_rsp_conv_51 = dat_rsp_conv_8b[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1562.4]
  assign dat_rsp_conv_52 = dat_rsp_conv_8b[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1564.4]
  assign dat_rsp_conv_53 = dat_rsp_conv_8b[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1566.4]
  assign dat_rsp_conv_54 = dat_rsp_conv_8b[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1568.4]
  assign dat_rsp_conv_55 = dat_rsp_conv_8b[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1570.4]
  assign dat_rsp_conv_56 = dat_rsp_conv_8b[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1572.4]
  assign dat_rsp_conv_57 = dat_rsp_conv_8b[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1574.4]
  assign dat_rsp_conv_58 = dat_rsp_conv_8b[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1576.4]
  assign dat_rsp_conv_59 = dat_rsp_conv_8b[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1578.4]
  assign dat_rsp_conv_60 = dat_rsp_conv_8b[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1580.4]
  assign dat_rsp_conv_61 = dat_rsp_conv_8b[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1582.4]
  assign dat_rsp_conv_62 = dat_rsp_conv_8b[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1584.4]
  assign dat_rsp_conv_63 = dat_rsp_conv_8b[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1057:39:@1586.4]
  assign _T_1834 = is_img_d1[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:39:@1594.4]
  assign _T_1835 = ~ _T_1834; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:29:@1595.4]
  assign _T_1837 = {dat_rsp_l0c0,dat_rsp_l0c1}; // @[Cat.scala 30:58:@1596.4]
  assign dat_rsp_l0_sft_in = _T_1835 ? 1024'h0 : _T_1837; // @[NV_NVDLA_CSC_dl_for_check.scala 1070:28:@1597.4]
  assign _T_1838 = is_img_d1[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1071:39:@1598.4]
  assign _T_1839 = ~ _T_1838; // @[NV_NVDLA_CSC_dl_for_check.scala 1071:29:@1599.4]
  assign _T_1841 = {dat_rsp_l1c0,dat_rsp_l1c1}; // @[Cat.scala 30:58:@1600.4]
  assign dat_rsp_l1_sft_in = _T_1839 ? 1024'h0 : _T_1841; // @[NV_NVDLA_CSC_dl_for_check.scala 1071:28:@1601.4]
  assign _T_1842 = is_img_d1[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:39:@1602.4]
  assign _T_1843 = ~ _T_1842; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:29:@1603.4]
  assign _T_1845 = {dat_rsp_l2c0,dat_rsp_l2c1}; // @[Cat.scala 30:58:@1604.4]
  assign dat_rsp_l2_sft_in = _T_1843 ? 1024'h0 : _T_1845; // @[NV_NVDLA_CSC_dl_for_check.scala 1072:28:@1605.4]
  assign _T_1846 = is_img_d1[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:39:@1606.4]
  assign _T_1847 = ~ _T_1846; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:29:@1607.4]
  assign _T_1849 = {dat_rsp_l3c0,dat_rsp_l3c1}; // @[Cat.scala 30:58:@1608.4]
  assign dat_rsp_l3_sft_in = _T_1847 ? 1024'h0 : _T_1849; // @[NV_NVDLA_CSC_dl_for_check.scala 1073:28:@1609.4]
  assign _T_1851 = {rsp_sft_cnt_l0,3'h0}; // @[Cat.scala 30:58:@1610.4]
  assign _T_1852 = dat_rsp_l0_sft_in >> _T_1851; // @[NV_NVDLA_CSC_dl_for_check.scala 1075:41:@1611.4]
  assign dat_rsp_l0_sft = _T_1852[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1075:82:@1612.4]
  assign _T_1854 = {rsp_sft_cnt_l1,3'h0}; // @[Cat.scala 30:58:@1613.4]
  assign _T_1855 = dat_rsp_l1_sft_in >> _T_1854; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:41:@1614.4]
  assign dat_rsp_l1_sft = _T_1855[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1076:82:@1615.4]
  assign _T_1857 = {rsp_sft_cnt_l2,3'h0}; // @[Cat.scala 30:58:@1616.4]
  assign _T_1858 = dat_rsp_l2_sft_in >> _T_1857; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:41:@1617.4]
  assign dat_rsp_l2_sft = _T_1858[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1077:82:@1618.4]
  assign _T_1860 = {rsp_sft_cnt_l3,3'h0}; // @[Cat.scala 30:58:@1619.4]
  assign _T_1861 = dat_rsp_l3_sft_in >> _T_1860; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:41:@1620.4]
  assign dat_rsp_l3_sft = _T_1861[511:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1078:82:@1621.4]
  assign _T_1862 = is_img_d1[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:36:@1622.4]
  assign _T_1863 = ~ _T_1862; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:26:@1623.4]
  assign _T_1866 = sub_h_total_g8 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1081:41:@1624.4]
  assign _T_1867 = dat_rsp_l3_sft[127:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1081:81:@1625.4]
  assign _T_1873 = {_T_1867,dat_rsp_l2_sft_d3,dat_rsp_l1_sft_d3,dat_rsp_l0_sft_d3}; // @[Cat.scala 30:58:@1631.4]
  assign _T_1875 = sub_h_total_g8 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:41:@1632.4]
  assign _T_1876 = dat_rsp_l1_sft[255:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:81:@1633.4]
  assign _T_1878 = {_T_1876,dat_rsp_l0_sft_d1}; // @[Cat.scala 30:58:@1635.4]
  assign _T_1880 = _T_1875 ? _T_1878 : dat_rsp_l0_sft; // @[NV_NVDLA_CSC_dl_for_check.scala 1082:25:@1637.4]
  assign _T_1881 = _T_1866 ? _T_1873 : _T_1880; // @[NV_NVDLA_CSC_dl_for_check.scala 1081:25:@1638.4]
  assign dat_rsp_img_8b = _T_1863 ? 512'h0 : _T_1881; // @[NV_NVDLA_CSC_dl_for_check.scala 1080:25:@1639.4]
  assign dat_rsp_img_0 = dat_rsp_img_8b[7:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1641.4]
  assign dat_rsp_img_1 = dat_rsp_img_8b[15:8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1643.4]
  assign dat_rsp_img_2 = dat_rsp_img_8b[23:16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1645.4]
  assign dat_rsp_img_3 = dat_rsp_img_8b[31:24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1647.4]
  assign dat_rsp_img_4 = dat_rsp_img_8b[39:32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1649.4]
  assign dat_rsp_img_5 = dat_rsp_img_8b[47:40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1651.4]
  assign dat_rsp_img_6 = dat_rsp_img_8b[55:48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1653.4]
  assign dat_rsp_img_7 = dat_rsp_img_8b[63:56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1655.4]
  assign dat_rsp_img_8 = dat_rsp_img_8b[71:64]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1657.4]
  assign dat_rsp_img_9 = dat_rsp_img_8b[79:72]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1659.4]
  assign dat_rsp_img_10 = dat_rsp_img_8b[87:80]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1661.4]
  assign dat_rsp_img_11 = dat_rsp_img_8b[95:88]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1663.4]
  assign dat_rsp_img_12 = dat_rsp_img_8b[103:96]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1665.4]
  assign dat_rsp_img_13 = dat_rsp_img_8b[111:104]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1667.4]
  assign dat_rsp_img_14 = dat_rsp_img_8b[119:112]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1669.4]
  assign dat_rsp_img_15 = dat_rsp_img_8b[127:120]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1671.4]
  assign dat_rsp_img_16 = dat_rsp_img_8b[135:128]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1673.4]
  assign dat_rsp_img_17 = dat_rsp_img_8b[143:136]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1675.4]
  assign dat_rsp_img_18 = dat_rsp_img_8b[151:144]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1677.4]
  assign dat_rsp_img_19 = dat_rsp_img_8b[159:152]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1679.4]
  assign dat_rsp_img_20 = dat_rsp_img_8b[167:160]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1681.4]
  assign dat_rsp_img_21 = dat_rsp_img_8b[175:168]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1683.4]
  assign dat_rsp_img_22 = dat_rsp_img_8b[183:176]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1685.4]
  assign dat_rsp_img_23 = dat_rsp_img_8b[191:184]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1687.4]
  assign dat_rsp_img_24 = dat_rsp_img_8b[199:192]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1689.4]
  assign dat_rsp_img_25 = dat_rsp_img_8b[207:200]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1691.4]
  assign dat_rsp_img_26 = dat_rsp_img_8b[215:208]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1693.4]
  assign dat_rsp_img_27 = dat_rsp_img_8b[223:216]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1695.4]
  assign dat_rsp_img_28 = dat_rsp_img_8b[231:224]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1697.4]
  assign dat_rsp_img_29 = dat_rsp_img_8b[239:232]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1699.4]
  assign dat_rsp_img_30 = dat_rsp_img_8b[247:240]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1701.4]
  assign dat_rsp_img_31 = dat_rsp_img_8b[255:248]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1703.4]
  assign dat_rsp_img_32 = dat_rsp_img_8b[263:256]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1705.4]
  assign dat_rsp_img_33 = dat_rsp_img_8b[271:264]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1707.4]
  assign dat_rsp_img_34 = dat_rsp_img_8b[279:272]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1709.4]
  assign dat_rsp_img_35 = dat_rsp_img_8b[287:280]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1711.4]
  assign dat_rsp_img_36 = dat_rsp_img_8b[295:288]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1713.4]
  assign dat_rsp_img_37 = dat_rsp_img_8b[303:296]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1715.4]
  assign dat_rsp_img_38 = dat_rsp_img_8b[311:304]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1717.4]
  assign dat_rsp_img_39 = dat_rsp_img_8b[319:312]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1719.4]
  assign dat_rsp_img_40 = dat_rsp_img_8b[327:320]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1721.4]
  assign dat_rsp_img_41 = dat_rsp_img_8b[335:328]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1723.4]
  assign dat_rsp_img_42 = dat_rsp_img_8b[343:336]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1725.4]
  assign dat_rsp_img_43 = dat_rsp_img_8b[351:344]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1727.4]
  assign dat_rsp_img_44 = dat_rsp_img_8b[359:352]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1729.4]
  assign dat_rsp_img_45 = dat_rsp_img_8b[367:360]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1731.4]
  assign dat_rsp_img_46 = dat_rsp_img_8b[375:368]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1733.4]
  assign dat_rsp_img_47 = dat_rsp_img_8b[383:376]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1735.4]
  assign dat_rsp_img_48 = dat_rsp_img_8b[391:384]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1737.4]
  assign dat_rsp_img_49 = dat_rsp_img_8b[399:392]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1739.4]
  assign dat_rsp_img_50 = dat_rsp_img_8b[407:400]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1741.4]
  assign dat_rsp_img_51 = dat_rsp_img_8b[415:408]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1743.4]
  assign dat_rsp_img_52 = dat_rsp_img_8b[423:416]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1745.4]
  assign dat_rsp_img_53 = dat_rsp_img_8b[431:424]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1747.4]
  assign dat_rsp_img_54 = dat_rsp_img_8b[439:432]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1749.4]
  assign dat_rsp_img_55 = dat_rsp_img_8b[447:440]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1751.4]
  assign dat_rsp_img_56 = dat_rsp_img_8b[455:448]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1753.4]
  assign dat_rsp_img_57 = dat_rsp_img_8b[463:456]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1755.4]
  assign dat_rsp_img_58 = dat_rsp_img_8b[471:464]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1757.4]
  assign dat_rsp_img_59 = dat_rsp_img_8b[479:472]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1759.4]
  assign dat_rsp_img_60 = dat_rsp_img_8b[487:480]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1761.4]
  assign dat_rsp_img_61 = dat_rsp_img_8b[495:488]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1763.4]
  assign dat_rsp_img_62 = dat_rsp_img_8b[503:496]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1765.4]
  assign dat_rsp_img_63 = dat_rsp_img_8b[511:504]; // @[NV_NVDLA_CSC_dl_for_check.scala 1088:37:@1767.4]
  assign _T_2016 = sub_h_total_g9 != 3'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1091:59:@1769.4]
  assign dat_rsp_sft_d1_en = dat_rsp_l0_pvld & _T_2016; // @[NV_NVDLA_CSC_dl_for_check.scala 1091:41:@1770.4]
  assign _T_2018 = sub_h_total_g9 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1092:59:@1771.4]
  assign dat_rsp_sft_d2_en = dat_rsp_l1_pvld & _T_2018; // @[NV_NVDLA_CSC_dl_for_check.scala 1092:41:@1772.4]
  assign dat_rsp_sft_d3_en = dat_rsp_l2_pvld & _T_2018; // @[NV_NVDLA_CSC_dl_for_check.scala 1093:41:@1774.4]
  assign _GEN_154 = dat_rsp_sft_d1_en ? dat_rsp_l0_sft : {{256'd0}, dat_rsp_l0_sft_d1}; // @[NV_NVDLA_CSC_dl_for_check.scala 1095:24:@1775.4]
  assign _GEN_155 = dat_rsp_sft_d2_en ? dat_rsp_l0_sft_d1 : {{128'd0}, dat_rsp_l0_sft_d2}; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:24:@1778.4]
  assign _GEN_156 = dat_rsp_sft_d2_en ? dat_rsp_l1_sft : {{384'd0}, dat_rsp_l1_sft_d2}; // @[NV_NVDLA_CSC_dl_for_check.scala 1098:24:@1778.4]
  assign _GEN_159 = dat_rsp_sft_d3_en ? dat_rsp_l2_sft : {{384'd0}, dat_rsp_l2_sft_d3}; // @[NV_NVDLA_CSC_dl_for_check.scala 1102:24:@1782.4]
  assign _T_2026 = 319'hffffffffffffffff << dat_rsp_bytes; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:55:@1788.4]
  assign dat_rsp_ori_mask = ~ _T_2026; // @[NV_NVDLA_CSC_dl_for_check.scala 1111:24:@1789.4]
  assign _T_2028 = dat_rsp_cur_sub_h >= 2'h1; // @[NV_NVDLA_CSC_dl_for_check.scala 1113:51:@1790.4]
  assign dat_rsp_cur_h_mask_p1 = _T_2028 ? 64'hffffffffffffffff : 64'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1113:32:@1792.4]
  assign _T_2036 = dat_rsp_cur_sub_h >= 2'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1114:51:@1793.4]
  assign dat_rsp_cur_h_mask_p2 = _T_2036 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1114:32:@1795.4]
  assign _T_2044 = dat_rsp_cur_sub_h == 2'h3; // @[NV_NVDLA_CSC_dl_for_check.scala 1115:51:@1796.4]
  assign dat_rsp_cur_h_mask_p3 = _T_2044 ? 32'hffffffff : 32'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1115:32:@1798.4]
  assign _T_2051 = dat_rsp_cur_h_mask_p1[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1117:57:@1799.4]
  assign dat_rsp_cur_h_e2_mask_8b = {_T_2051,32'hffffffff}; // @[Cat.scala 30:58:@1801.4]
  assign _T_2057 = dat_rsp_cur_h_mask_p3[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:57:@1802.4]
  assign _T_2058 = dat_rsp_cur_h_mask_p2[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:106:@1803.4]
  assign _T_2059 = dat_rsp_cur_h_mask_p1[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1118:155:@1804.4]
  assign dat_rsp_cur_h_e4_mask_8b = {_T_2057,_T_2058,_T_2059,16'hffff}; // @[Cat.scala 30:58:@1808.4]
  assign _T_2068 = sub_h_total_g11 == 3'h4; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:43:@1809.4]
  assign _T_2069 = dat_rsp_ori_mask[15:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:89:@1810.4]
  assign _T_2071 = {_T_2069,_T_2069,_T_2069,_T_2069}; // @[Cat.scala 30:58:@1812.4]
  assign _T_2072 = _T_2071 & dat_rsp_cur_h_e4_mask_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:116:@1813.4]
  assign _T_2074 = sub_h_total_g11 == 3'h2; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:43:@1814.4]
  assign _T_2075 = dat_rsp_ori_mask[31:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:89:@1815.4]
  assign _T_2076 = {_T_2075,_T_2075}; // @[Cat.scala 30:58:@1816.4]
  assign _T_2077 = _T_2076 & dat_rsp_cur_h_e2_mask_8b; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:116:@1817.4]
  assign _T_2078 = dat_rsp_ori_mask[63:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1122:39:@1818.4]
  assign _T_2079 = _T_2074 ? _T_2077 : _T_2078; // @[NV_NVDLA_CSC_dl_for_check.scala 1121:26:@1819.4]
  assign dat_rsp_mask_8b = _T_2068 ? _T_2072 : _T_2079; // @[NV_NVDLA_CSC_dl_for_check.scala 1120:26:@1820.4]
  assign _T_2080 = is_img_d1[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:35:@1821.4]
  assign dat_rsp_data_w_0 = _T_2080 ? dat_rsp_img_0 : dat_rsp_conv_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_1 = _T_2080 ? dat_rsp_img_1 : dat_rsp_conv_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_2 = _T_2080 ? dat_rsp_img_2 : dat_rsp_conv_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_3 = _T_2080 ? dat_rsp_img_3 : dat_rsp_conv_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_4 = _T_2080 ? dat_rsp_img_4 : dat_rsp_conv_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_5 = _T_2080 ? dat_rsp_img_5 : dat_rsp_conv_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_6 = _T_2080 ? dat_rsp_img_6 : dat_rsp_conv_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_7 = _T_2080 ? dat_rsp_img_7 : dat_rsp_conv_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_8 = _T_2080 ? dat_rsp_img_8 : dat_rsp_conv_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_9 = _T_2080 ? dat_rsp_img_9 : dat_rsp_conv_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_10 = _T_2080 ? dat_rsp_img_10 : dat_rsp_conv_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_11 = _T_2080 ? dat_rsp_img_11 : dat_rsp_conv_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_12 = _T_2080 ? dat_rsp_img_12 : dat_rsp_conv_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_13 = _T_2080 ? dat_rsp_img_13 : dat_rsp_conv_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_14 = _T_2080 ? dat_rsp_img_14 : dat_rsp_conv_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_15 = _T_2080 ? dat_rsp_img_15 : dat_rsp_conv_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_16 = _T_2080 ? dat_rsp_img_16 : dat_rsp_conv_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_17 = _T_2080 ? dat_rsp_img_17 : dat_rsp_conv_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_18 = _T_2080 ? dat_rsp_img_18 : dat_rsp_conv_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_19 = _T_2080 ? dat_rsp_img_19 : dat_rsp_conv_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_20 = _T_2080 ? dat_rsp_img_20 : dat_rsp_conv_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_21 = _T_2080 ? dat_rsp_img_21 : dat_rsp_conv_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_22 = _T_2080 ? dat_rsp_img_22 : dat_rsp_conv_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_23 = _T_2080 ? dat_rsp_img_23 : dat_rsp_conv_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_24 = _T_2080 ? dat_rsp_img_24 : dat_rsp_conv_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_25 = _T_2080 ? dat_rsp_img_25 : dat_rsp_conv_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_26 = _T_2080 ? dat_rsp_img_26 : dat_rsp_conv_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_27 = _T_2080 ? dat_rsp_img_27 : dat_rsp_conv_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_28 = _T_2080 ? dat_rsp_img_28 : dat_rsp_conv_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_29 = _T_2080 ? dat_rsp_img_29 : dat_rsp_conv_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_30 = _T_2080 ? dat_rsp_img_30 : dat_rsp_conv_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_31 = _T_2080 ? dat_rsp_img_31 : dat_rsp_conv_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_32 = _T_2080 ? dat_rsp_img_32 : dat_rsp_conv_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_33 = _T_2080 ? dat_rsp_img_33 : dat_rsp_conv_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_34 = _T_2080 ? dat_rsp_img_34 : dat_rsp_conv_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_35 = _T_2080 ? dat_rsp_img_35 : dat_rsp_conv_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_36 = _T_2080 ? dat_rsp_img_36 : dat_rsp_conv_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_37 = _T_2080 ? dat_rsp_img_37 : dat_rsp_conv_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_38 = _T_2080 ? dat_rsp_img_38 : dat_rsp_conv_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_39 = _T_2080 ? dat_rsp_img_39 : dat_rsp_conv_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_40 = _T_2080 ? dat_rsp_img_40 : dat_rsp_conv_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_41 = _T_2080 ? dat_rsp_img_41 : dat_rsp_conv_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_42 = _T_2080 ? dat_rsp_img_42 : dat_rsp_conv_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_43 = _T_2080 ? dat_rsp_img_43 : dat_rsp_conv_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_44 = _T_2080 ? dat_rsp_img_44 : dat_rsp_conv_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_45 = _T_2080 ? dat_rsp_img_45 : dat_rsp_conv_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_46 = _T_2080 ? dat_rsp_img_46 : dat_rsp_conv_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_47 = _T_2080 ? dat_rsp_img_47 : dat_rsp_conv_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_48 = _T_2080 ? dat_rsp_img_48 : dat_rsp_conv_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_49 = _T_2080 ? dat_rsp_img_49 : dat_rsp_conv_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_50 = _T_2080 ? dat_rsp_img_50 : dat_rsp_conv_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_51 = _T_2080 ? dat_rsp_img_51 : dat_rsp_conv_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_52 = _T_2080 ? dat_rsp_img_52 : dat_rsp_conv_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_53 = _T_2080 ? dat_rsp_img_53 : dat_rsp_conv_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_54 = _T_2080 ? dat_rsp_img_54 : dat_rsp_conv_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_55 = _T_2080 ? dat_rsp_img_55 : dat_rsp_conv_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_56 = _T_2080 ? dat_rsp_img_56 : dat_rsp_conv_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_57 = _T_2080 ? dat_rsp_img_57 : dat_rsp_conv_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_58 = _T_2080 ? dat_rsp_img_58 : dat_rsp_conv_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_59 = _T_2080 ? dat_rsp_img_59 : dat_rsp_conv_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_60 = _T_2080 ? dat_rsp_img_60 : dat_rsp_conv_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_61 = _T_2080 ? dat_rsp_img_61 : dat_rsp_conv_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_62 = _T_2080 ? dat_rsp_img_62 : dat_rsp_conv_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_data_w_63 = _T_2080 ? dat_rsp_img_63 : dat_rsp_conv_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1125:25:@1822.4]
  assign dat_rsp_mask_val_int8_0 = dat_rsp_data_w_0 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1823.4]
  assign dat_rsp_mask_val_int8_1 = dat_rsp_data_w_1 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1824.4]
  assign dat_rsp_mask_val_int8_2 = dat_rsp_data_w_2 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1825.4]
  assign dat_rsp_mask_val_int8_3 = dat_rsp_data_w_3 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1826.4]
  assign dat_rsp_mask_val_int8_4 = dat_rsp_data_w_4 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1827.4]
  assign dat_rsp_mask_val_int8_5 = dat_rsp_data_w_5 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1828.4]
  assign dat_rsp_mask_val_int8_6 = dat_rsp_data_w_6 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1829.4]
  assign dat_rsp_mask_val_int8_7 = dat_rsp_data_w_7 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1830.4]
  assign dat_rsp_mask_val_int8_8 = dat_rsp_data_w_8 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1831.4]
  assign dat_rsp_mask_val_int8_9 = dat_rsp_data_w_9 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1832.4]
  assign dat_rsp_mask_val_int8_10 = dat_rsp_data_w_10 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1833.4]
  assign dat_rsp_mask_val_int8_11 = dat_rsp_data_w_11 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1834.4]
  assign dat_rsp_mask_val_int8_12 = dat_rsp_data_w_12 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1835.4]
  assign dat_rsp_mask_val_int8_13 = dat_rsp_data_w_13 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1836.4]
  assign dat_rsp_mask_val_int8_14 = dat_rsp_data_w_14 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1837.4]
  assign dat_rsp_mask_val_int8_15 = dat_rsp_data_w_15 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1838.4]
  assign dat_rsp_mask_val_int8_16 = dat_rsp_data_w_16 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1839.4]
  assign dat_rsp_mask_val_int8_17 = dat_rsp_data_w_17 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1840.4]
  assign dat_rsp_mask_val_int8_18 = dat_rsp_data_w_18 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1841.4]
  assign dat_rsp_mask_val_int8_19 = dat_rsp_data_w_19 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1842.4]
  assign dat_rsp_mask_val_int8_20 = dat_rsp_data_w_20 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1843.4]
  assign dat_rsp_mask_val_int8_21 = dat_rsp_data_w_21 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1844.4]
  assign dat_rsp_mask_val_int8_22 = dat_rsp_data_w_22 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1845.4]
  assign dat_rsp_mask_val_int8_23 = dat_rsp_data_w_23 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1846.4]
  assign dat_rsp_mask_val_int8_24 = dat_rsp_data_w_24 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1847.4]
  assign dat_rsp_mask_val_int8_25 = dat_rsp_data_w_25 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1848.4]
  assign dat_rsp_mask_val_int8_26 = dat_rsp_data_w_26 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1849.4]
  assign dat_rsp_mask_val_int8_27 = dat_rsp_data_w_27 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1850.4]
  assign dat_rsp_mask_val_int8_28 = dat_rsp_data_w_28 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1851.4]
  assign dat_rsp_mask_val_int8_29 = dat_rsp_data_w_29 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1852.4]
  assign dat_rsp_mask_val_int8_30 = dat_rsp_data_w_30 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1853.4]
  assign dat_rsp_mask_val_int8_31 = dat_rsp_data_w_31 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1854.4]
  assign dat_rsp_mask_val_int8_32 = dat_rsp_data_w_32 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1855.4]
  assign dat_rsp_mask_val_int8_33 = dat_rsp_data_w_33 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1856.4]
  assign dat_rsp_mask_val_int8_34 = dat_rsp_data_w_34 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1857.4]
  assign dat_rsp_mask_val_int8_35 = dat_rsp_data_w_35 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1858.4]
  assign dat_rsp_mask_val_int8_36 = dat_rsp_data_w_36 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1859.4]
  assign dat_rsp_mask_val_int8_37 = dat_rsp_data_w_37 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1860.4]
  assign dat_rsp_mask_val_int8_38 = dat_rsp_data_w_38 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1861.4]
  assign dat_rsp_mask_val_int8_39 = dat_rsp_data_w_39 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1862.4]
  assign dat_rsp_mask_val_int8_40 = dat_rsp_data_w_40 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1863.4]
  assign dat_rsp_mask_val_int8_41 = dat_rsp_data_w_41 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1864.4]
  assign dat_rsp_mask_val_int8_42 = dat_rsp_data_w_42 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1865.4]
  assign dat_rsp_mask_val_int8_43 = dat_rsp_data_w_43 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1866.4]
  assign dat_rsp_mask_val_int8_44 = dat_rsp_data_w_44 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1867.4]
  assign dat_rsp_mask_val_int8_45 = dat_rsp_data_w_45 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1868.4]
  assign dat_rsp_mask_val_int8_46 = dat_rsp_data_w_46 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1869.4]
  assign dat_rsp_mask_val_int8_47 = dat_rsp_data_w_47 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1870.4]
  assign dat_rsp_mask_val_int8_48 = dat_rsp_data_w_48 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1871.4]
  assign dat_rsp_mask_val_int8_49 = dat_rsp_data_w_49 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1872.4]
  assign dat_rsp_mask_val_int8_50 = dat_rsp_data_w_50 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1873.4]
  assign dat_rsp_mask_val_int8_51 = dat_rsp_data_w_51 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1874.4]
  assign dat_rsp_mask_val_int8_52 = dat_rsp_data_w_52 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1875.4]
  assign dat_rsp_mask_val_int8_53 = dat_rsp_data_w_53 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1876.4]
  assign dat_rsp_mask_val_int8_54 = dat_rsp_data_w_54 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1877.4]
  assign dat_rsp_mask_val_int8_55 = dat_rsp_data_w_55 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1878.4]
  assign dat_rsp_mask_val_int8_56 = dat_rsp_data_w_56 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1879.4]
  assign dat_rsp_mask_val_int8_57 = dat_rsp_data_w_57 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1880.4]
  assign dat_rsp_mask_val_int8_58 = dat_rsp_data_w_58 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1881.4]
  assign dat_rsp_mask_val_int8_59 = dat_rsp_data_w_59 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1882.4]
  assign dat_rsp_mask_val_int8_60 = dat_rsp_data_w_60 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1883.4]
  assign dat_rsp_mask_val_int8_61 = dat_rsp_data_w_61 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1884.4]
  assign dat_rsp_mask_val_int8_62 = dat_rsp_data_w_62 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1885.4]
  assign dat_rsp_mask_val_int8_63 = dat_rsp_data_w_63 != 8'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 1126:97:@1886.4]
  assign _T_2409 = dat_rsp_mask_8b[0]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1952.4]
  assign dat_rsp_mask_w_0 = _T_2409 & dat_rsp_mask_val_int8_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1953.4]
  assign _T_2411 = dat_rsp_mask_8b[1]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1954.4]
  assign dat_rsp_mask_w_1 = _T_2411 & dat_rsp_mask_val_int8_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1955.4]
  assign _T_2413 = dat_rsp_mask_8b[2]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1956.4]
  assign dat_rsp_mask_w_2 = _T_2413 & dat_rsp_mask_val_int8_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1957.4]
  assign _T_2415 = dat_rsp_mask_8b[3]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1958.4]
  assign dat_rsp_mask_w_3 = _T_2415 & dat_rsp_mask_val_int8_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1959.4]
  assign _T_2417 = dat_rsp_mask_8b[4]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1960.4]
  assign dat_rsp_mask_w_4 = _T_2417 & dat_rsp_mask_val_int8_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1961.4]
  assign _T_2419 = dat_rsp_mask_8b[5]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1962.4]
  assign dat_rsp_mask_w_5 = _T_2419 & dat_rsp_mask_val_int8_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1963.4]
  assign _T_2421 = dat_rsp_mask_8b[6]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1964.4]
  assign dat_rsp_mask_w_6 = _T_2421 & dat_rsp_mask_val_int8_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1965.4]
  assign _T_2423 = dat_rsp_mask_8b[7]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1966.4]
  assign dat_rsp_mask_w_7 = _T_2423 & dat_rsp_mask_val_int8_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1967.4]
  assign _T_2425 = dat_rsp_mask_8b[8]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1968.4]
  assign dat_rsp_mask_w_8 = _T_2425 & dat_rsp_mask_val_int8_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1969.4]
  assign _T_2427 = dat_rsp_mask_8b[9]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1970.4]
  assign dat_rsp_mask_w_9 = _T_2427 & dat_rsp_mask_val_int8_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1971.4]
  assign _T_2429 = dat_rsp_mask_8b[10]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1972.4]
  assign dat_rsp_mask_w_10 = _T_2429 & dat_rsp_mask_val_int8_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1973.4]
  assign _T_2431 = dat_rsp_mask_8b[11]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1974.4]
  assign dat_rsp_mask_w_11 = _T_2431 & dat_rsp_mask_val_int8_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1975.4]
  assign _T_2433 = dat_rsp_mask_8b[12]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1976.4]
  assign dat_rsp_mask_w_12 = _T_2433 & dat_rsp_mask_val_int8_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1977.4]
  assign _T_2435 = dat_rsp_mask_8b[13]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1978.4]
  assign dat_rsp_mask_w_13 = _T_2435 & dat_rsp_mask_val_int8_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1979.4]
  assign _T_2437 = dat_rsp_mask_8b[14]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1980.4]
  assign dat_rsp_mask_w_14 = _T_2437 & dat_rsp_mask_val_int8_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1981.4]
  assign _T_2439 = dat_rsp_mask_8b[15]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1982.4]
  assign dat_rsp_mask_w_15 = _T_2439 & dat_rsp_mask_val_int8_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1983.4]
  assign _T_2441 = dat_rsp_mask_8b[16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1984.4]
  assign dat_rsp_mask_w_16 = _T_2441 & dat_rsp_mask_val_int8_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1985.4]
  assign _T_2443 = dat_rsp_mask_8b[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1986.4]
  assign dat_rsp_mask_w_17 = _T_2443 & dat_rsp_mask_val_int8_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1987.4]
  assign _T_2445 = dat_rsp_mask_8b[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1988.4]
  assign dat_rsp_mask_w_18 = _T_2445 & dat_rsp_mask_val_int8_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1989.4]
  assign _T_2447 = dat_rsp_mask_8b[19]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1990.4]
  assign dat_rsp_mask_w_19 = _T_2447 & dat_rsp_mask_val_int8_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1991.4]
  assign _T_2449 = dat_rsp_mask_8b[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1992.4]
  assign dat_rsp_mask_w_20 = _T_2449 & dat_rsp_mask_val_int8_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1993.4]
  assign _T_2451 = dat_rsp_mask_8b[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1994.4]
  assign dat_rsp_mask_w_21 = _T_2451 & dat_rsp_mask_val_int8_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1995.4]
  assign _T_2453 = dat_rsp_mask_8b[22]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1996.4]
  assign dat_rsp_mask_w_22 = _T_2453 & dat_rsp_mask_val_int8_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1997.4]
  assign _T_2455 = dat_rsp_mask_8b[23]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@1998.4]
  assign dat_rsp_mask_w_23 = _T_2455 & dat_rsp_mask_val_int8_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@1999.4]
  assign _T_2457 = dat_rsp_mask_8b[24]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2000.4]
  assign dat_rsp_mask_w_24 = _T_2457 & dat_rsp_mask_val_int8_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2001.4]
  assign _T_2459 = dat_rsp_mask_8b[25]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2002.4]
  assign dat_rsp_mask_w_25 = _T_2459 & dat_rsp_mask_val_int8_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2003.4]
  assign _T_2461 = dat_rsp_mask_8b[26]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2004.4]
  assign dat_rsp_mask_w_26 = _T_2461 & dat_rsp_mask_val_int8_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2005.4]
  assign _T_2463 = dat_rsp_mask_8b[27]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2006.4]
  assign dat_rsp_mask_w_27 = _T_2463 & dat_rsp_mask_val_int8_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2007.4]
  assign _T_2465 = dat_rsp_mask_8b[28]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2008.4]
  assign dat_rsp_mask_w_28 = _T_2465 & dat_rsp_mask_val_int8_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2009.4]
  assign _T_2467 = dat_rsp_mask_8b[29]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2010.4]
  assign dat_rsp_mask_w_29 = _T_2467 & dat_rsp_mask_val_int8_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2011.4]
  assign _T_2469 = dat_rsp_mask_8b[30]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2012.4]
  assign dat_rsp_mask_w_30 = _T_2469 & dat_rsp_mask_val_int8_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2013.4]
  assign _T_2471 = dat_rsp_mask_8b[31]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2014.4]
  assign dat_rsp_mask_w_31 = _T_2471 & dat_rsp_mask_val_int8_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2015.4]
  assign _T_2473 = dat_rsp_mask_8b[32]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2016.4]
  assign dat_rsp_mask_w_32 = _T_2473 & dat_rsp_mask_val_int8_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2017.4]
  assign _T_2475 = dat_rsp_mask_8b[33]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2018.4]
  assign dat_rsp_mask_w_33 = _T_2475 & dat_rsp_mask_val_int8_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2019.4]
  assign _T_2477 = dat_rsp_mask_8b[34]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2020.4]
  assign dat_rsp_mask_w_34 = _T_2477 & dat_rsp_mask_val_int8_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2021.4]
  assign _T_2479 = dat_rsp_mask_8b[35]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2022.4]
  assign dat_rsp_mask_w_35 = _T_2479 & dat_rsp_mask_val_int8_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2023.4]
  assign _T_2481 = dat_rsp_mask_8b[36]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2024.4]
  assign dat_rsp_mask_w_36 = _T_2481 & dat_rsp_mask_val_int8_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2025.4]
  assign _T_2483 = dat_rsp_mask_8b[37]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2026.4]
  assign dat_rsp_mask_w_37 = _T_2483 & dat_rsp_mask_val_int8_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2027.4]
  assign _T_2485 = dat_rsp_mask_8b[38]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2028.4]
  assign dat_rsp_mask_w_38 = _T_2485 & dat_rsp_mask_val_int8_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2029.4]
  assign _T_2487 = dat_rsp_mask_8b[39]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2030.4]
  assign dat_rsp_mask_w_39 = _T_2487 & dat_rsp_mask_val_int8_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2031.4]
  assign _T_2489 = dat_rsp_mask_8b[40]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2032.4]
  assign dat_rsp_mask_w_40 = _T_2489 & dat_rsp_mask_val_int8_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2033.4]
  assign _T_2491 = dat_rsp_mask_8b[41]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2034.4]
  assign dat_rsp_mask_w_41 = _T_2491 & dat_rsp_mask_val_int8_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2035.4]
  assign _T_2493 = dat_rsp_mask_8b[42]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2036.4]
  assign dat_rsp_mask_w_42 = _T_2493 & dat_rsp_mask_val_int8_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2037.4]
  assign _T_2495 = dat_rsp_mask_8b[43]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2038.4]
  assign dat_rsp_mask_w_43 = _T_2495 & dat_rsp_mask_val_int8_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2039.4]
  assign _T_2497 = dat_rsp_mask_8b[44]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2040.4]
  assign dat_rsp_mask_w_44 = _T_2497 & dat_rsp_mask_val_int8_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2041.4]
  assign _T_2499 = dat_rsp_mask_8b[45]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2042.4]
  assign dat_rsp_mask_w_45 = _T_2499 & dat_rsp_mask_val_int8_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2043.4]
  assign _T_2501 = dat_rsp_mask_8b[46]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2044.4]
  assign dat_rsp_mask_w_46 = _T_2501 & dat_rsp_mask_val_int8_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2045.4]
  assign _T_2503 = dat_rsp_mask_8b[47]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2046.4]
  assign dat_rsp_mask_w_47 = _T_2503 & dat_rsp_mask_val_int8_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2047.4]
  assign _T_2505 = dat_rsp_mask_8b[48]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2048.4]
  assign dat_rsp_mask_w_48 = _T_2505 & dat_rsp_mask_val_int8_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2049.4]
  assign _T_2507 = dat_rsp_mask_8b[49]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2050.4]
  assign dat_rsp_mask_w_49 = _T_2507 & dat_rsp_mask_val_int8_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2051.4]
  assign _T_2509 = dat_rsp_mask_8b[50]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2052.4]
  assign dat_rsp_mask_w_50 = _T_2509 & dat_rsp_mask_val_int8_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2053.4]
  assign _T_2511 = dat_rsp_mask_8b[51]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2054.4]
  assign dat_rsp_mask_w_51 = _T_2511 & dat_rsp_mask_val_int8_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2055.4]
  assign _T_2513 = dat_rsp_mask_8b[52]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2056.4]
  assign dat_rsp_mask_w_52 = _T_2513 & dat_rsp_mask_val_int8_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2057.4]
  assign _T_2515 = dat_rsp_mask_8b[53]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2058.4]
  assign dat_rsp_mask_w_53 = _T_2515 & dat_rsp_mask_val_int8_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2059.4]
  assign _T_2517 = dat_rsp_mask_8b[54]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2060.4]
  assign dat_rsp_mask_w_54 = _T_2517 & dat_rsp_mask_val_int8_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2061.4]
  assign _T_2519 = dat_rsp_mask_8b[55]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2062.4]
  assign dat_rsp_mask_w_55 = _T_2519 & dat_rsp_mask_val_int8_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2063.4]
  assign _T_2521 = dat_rsp_mask_8b[56]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2064.4]
  assign dat_rsp_mask_w_56 = _T_2521 & dat_rsp_mask_val_int8_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2065.4]
  assign _T_2523 = dat_rsp_mask_8b[57]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2066.4]
  assign dat_rsp_mask_w_57 = _T_2523 & dat_rsp_mask_val_int8_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2067.4]
  assign _T_2525 = dat_rsp_mask_8b[58]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2068.4]
  assign dat_rsp_mask_w_58 = _T_2525 & dat_rsp_mask_val_int8_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2069.4]
  assign _T_2527 = dat_rsp_mask_8b[59]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2070.4]
  assign dat_rsp_mask_w_59 = _T_2527 & dat_rsp_mask_val_int8_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2071.4]
  assign _T_2529 = dat_rsp_mask_8b[60]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2072.4]
  assign dat_rsp_mask_w_60 = _T_2529 & dat_rsp_mask_val_int8_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2073.4]
  assign _T_2531 = dat_rsp_mask_8b[61]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2074.4]
  assign dat_rsp_mask_w_61 = _T_2531 & dat_rsp_mask_val_int8_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2075.4]
  assign _T_2533 = dat_rsp_mask_8b[62]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2076.4]
  assign dat_rsp_mask_w_62 = _T_2533 & dat_rsp_mask_val_int8_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2077.4]
  assign _T_2535 = dat_rsp_mask_8b[63]; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:80:@2078.4]
  assign dat_rsp_mask_w_63 = _T_2535 & dat_rsp_mask_val_int8_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1127:83:@2079.4]
  assign _T_2606 = is_winograd_d1[16]; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:54:@2145.4]
  assign _T_2607 = ~ _T_2606; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:39:@2146.4]
  assign dat_rsp_p0_vld_w = dat_rsp_pvld & _T_2607; // @[NV_NVDLA_CSC_dl_for_check.scala 1128:37:@2147.4]
  assign _GEN_160 = dat_rsp_pvld ? dat_rsp_flag : _T_3164; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2232.4]
  assign _GEN_161 = _T_3147 ? _T_3164 : _T_3167; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2236.4]
  assign _GEN_162 = _T_3150 ? _T_3167 : _T_3170; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2240.4]
  assign _GEN_163 = _T_3153 ? _T_3170 : _T_3173; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2244.4]
  assign _GEN_164 = _T_3156 ? _T_3173 : _T_3176; // @[NV_NVDLA_CSC_dl_for_check.scala 1148:28:@2248.4]
  assign _T_3177 = is_winograd_d1[17]; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:40:@2251.4]
  assign dat_out_pvld_w = _T_3177 ? _T_3159 : dat_rsp_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1153:25:@2252.4]
  assign _T_3178 = is_winograd_d1[18]; // @[NV_NVDLA_CSC_dl_for_check.scala 1154:40:@2253.4]
  assign dat_out_flag_w = _T_3178 ? _T_3176 : dat_rsp_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1154:25:@2254.4]
  assign _GEN_165 = dat_out_pvld_w ? dat_out_flag_w : dat_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1161:21:@2256.4]
  assign _GEN_166 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_0 : dat_out_bypass_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_167 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_1 : dat_out_bypass_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_168 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_2 : dat_out_bypass_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_169 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_3 : dat_out_bypass_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_170 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_4 : dat_out_bypass_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_171 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_5 : dat_out_bypass_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_172 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_6 : dat_out_bypass_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_173 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_7 : dat_out_bypass_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_174 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_8 : dat_out_bypass_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_175 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_9 : dat_out_bypass_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_176 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_10 : dat_out_bypass_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_177 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_11 : dat_out_bypass_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_178 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_12 : dat_out_bypass_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_179 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_13 : dat_out_bypass_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_180 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_14 : dat_out_bypass_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_181 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_15 : dat_out_bypass_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_182 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_16 : dat_out_bypass_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_183 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_17 : dat_out_bypass_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_184 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_18 : dat_out_bypass_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_185 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_19 : dat_out_bypass_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_186 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_20 : dat_out_bypass_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_187 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_21 : dat_out_bypass_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_188 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_22 : dat_out_bypass_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_189 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_23 : dat_out_bypass_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_190 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_24 : dat_out_bypass_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_191 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_25 : dat_out_bypass_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_192 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_26 : dat_out_bypass_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_193 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_27 : dat_out_bypass_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_194 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_28 : dat_out_bypass_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_195 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_29 : dat_out_bypass_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_196 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_30 : dat_out_bypass_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_197 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_31 : dat_out_bypass_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_198 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_32 : dat_out_bypass_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_199 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_33 : dat_out_bypass_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_200 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_34 : dat_out_bypass_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_201 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_35 : dat_out_bypass_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_202 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_36 : dat_out_bypass_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_203 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_37 : dat_out_bypass_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_204 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_38 : dat_out_bypass_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_205 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_39 : dat_out_bypass_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_206 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_40 : dat_out_bypass_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_207 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_41 : dat_out_bypass_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_208 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_42 : dat_out_bypass_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_209 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_43 : dat_out_bypass_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_210 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_44 : dat_out_bypass_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_211 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_45 : dat_out_bypass_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_212 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_46 : dat_out_bypass_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_213 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_47 : dat_out_bypass_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_214 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_48 : dat_out_bypass_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_215 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_49 : dat_out_bypass_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_216 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_50 : dat_out_bypass_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_217 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_51 : dat_out_bypass_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_218 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_52 : dat_out_bypass_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_219 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_53 : dat_out_bypass_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_220 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_54 : dat_out_bypass_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_221 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_55 : dat_out_bypass_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_222 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_56 : dat_out_bypass_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_223 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_57 : dat_out_bypass_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_224 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_58 : dat_out_bypass_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_225 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_59 : dat_out_bypass_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_226 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_60 : dat_out_bypass_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_227 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_61 : dat_out_bypass_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_228 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_62 : dat_out_bypass_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _GEN_229 = dat_rsp_p0_vld_w ? dat_rsp_mask_w_63 : dat_out_bypass_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1164:30:@2259.4]
  assign _T_3179 = dat_rsp_p0_vld_w & dat_rsp_mask_w_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2325.4]
  assign _T_3180 = dat_rsp_p0_vld_w & dat_rsp_mask_w_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2329.4]
  assign _T_3181 = dat_rsp_p0_vld_w & dat_rsp_mask_w_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2333.4]
  assign _T_3182 = dat_rsp_p0_vld_w & dat_rsp_mask_w_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2337.4]
  assign _T_3183 = dat_rsp_p0_vld_w & dat_rsp_mask_w_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2341.4]
  assign _T_3184 = dat_rsp_p0_vld_w & dat_rsp_mask_w_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2345.4]
  assign _T_3185 = dat_rsp_p0_vld_w & dat_rsp_mask_w_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2349.4]
  assign _T_3186 = dat_rsp_p0_vld_w & dat_rsp_mask_w_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2353.4]
  assign _T_3187 = dat_rsp_p0_vld_w & dat_rsp_mask_w_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2357.4]
  assign _T_3188 = dat_rsp_p0_vld_w & dat_rsp_mask_w_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2361.4]
  assign _T_3189 = dat_rsp_p0_vld_w & dat_rsp_mask_w_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2365.4]
  assign _T_3190 = dat_rsp_p0_vld_w & dat_rsp_mask_w_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2369.4]
  assign _T_3191 = dat_rsp_p0_vld_w & dat_rsp_mask_w_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2373.4]
  assign _T_3192 = dat_rsp_p0_vld_w & dat_rsp_mask_w_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2377.4]
  assign _T_3193 = dat_rsp_p0_vld_w & dat_rsp_mask_w_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2381.4]
  assign _T_3194 = dat_rsp_p0_vld_w & dat_rsp_mask_w_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2385.4]
  assign _T_3195 = dat_rsp_p0_vld_w & dat_rsp_mask_w_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2389.4]
  assign _T_3196 = dat_rsp_p0_vld_w & dat_rsp_mask_w_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2393.4]
  assign _T_3197 = dat_rsp_p0_vld_w & dat_rsp_mask_w_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2397.4]
  assign _T_3198 = dat_rsp_p0_vld_w & dat_rsp_mask_w_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2401.4]
  assign _T_3199 = dat_rsp_p0_vld_w & dat_rsp_mask_w_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2405.4]
  assign _T_3200 = dat_rsp_p0_vld_w & dat_rsp_mask_w_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2409.4]
  assign _T_3201 = dat_rsp_p0_vld_w & dat_rsp_mask_w_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2413.4]
  assign _T_3202 = dat_rsp_p0_vld_w & dat_rsp_mask_w_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2417.4]
  assign _T_3203 = dat_rsp_p0_vld_w & dat_rsp_mask_w_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2421.4]
  assign _T_3204 = dat_rsp_p0_vld_w & dat_rsp_mask_w_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2425.4]
  assign _T_3205 = dat_rsp_p0_vld_w & dat_rsp_mask_w_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2429.4]
  assign _T_3206 = dat_rsp_p0_vld_w & dat_rsp_mask_w_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2433.4]
  assign _T_3207 = dat_rsp_p0_vld_w & dat_rsp_mask_w_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2437.4]
  assign _T_3208 = dat_rsp_p0_vld_w & dat_rsp_mask_w_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2441.4]
  assign _T_3209 = dat_rsp_p0_vld_w & dat_rsp_mask_w_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2445.4]
  assign _T_3210 = dat_rsp_p0_vld_w & dat_rsp_mask_w_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2449.4]
  assign _T_3211 = dat_rsp_p0_vld_w & dat_rsp_mask_w_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2453.4]
  assign _T_3212 = dat_rsp_p0_vld_w & dat_rsp_mask_w_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2457.4]
  assign _T_3213 = dat_rsp_p0_vld_w & dat_rsp_mask_w_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2461.4]
  assign _T_3214 = dat_rsp_p0_vld_w & dat_rsp_mask_w_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2465.4]
  assign _T_3215 = dat_rsp_p0_vld_w & dat_rsp_mask_w_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2469.4]
  assign _T_3216 = dat_rsp_p0_vld_w & dat_rsp_mask_w_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2473.4]
  assign _T_3217 = dat_rsp_p0_vld_w & dat_rsp_mask_w_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2477.4]
  assign _T_3218 = dat_rsp_p0_vld_w & dat_rsp_mask_w_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2481.4]
  assign _T_3219 = dat_rsp_p0_vld_w & dat_rsp_mask_w_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2485.4]
  assign _T_3220 = dat_rsp_p0_vld_w & dat_rsp_mask_w_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2489.4]
  assign _T_3221 = dat_rsp_p0_vld_w & dat_rsp_mask_w_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2493.4]
  assign _T_3222 = dat_rsp_p0_vld_w & dat_rsp_mask_w_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2497.4]
  assign _T_3223 = dat_rsp_p0_vld_w & dat_rsp_mask_w_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2501.4]
  assign _T_3224 = dat_rsp_p0_vld_w & dat_rsp_mask_w_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2505.4]
  assign _T_3225 = dat_rsp_p0_vld_w & dat_rsp_mask_w_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2509.4]
  assign _T_3226 = dat_rsp_p0_vld_w & dat_rsp_mask_w_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2513.4]
  assign _T_3227 = dat_rsp_p0_vld_w & dat_rsp_mask_w_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2517.4]
  assign _T_3228 = dat_rsp_p0_vld_w & dat_rsp_mask_w_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2521.4]
  assign _T_3229 = dat_rsp_p0_vld_w & dat_rsp_mask_w_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2525.4]
  assign _T_3230 = dat_rsp_p0_vld_w & dat_rsp_mask_w_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2529.4]
  assign _T_3231 = dat_rsp_p0_vld_w & dat_rsp_mask_w_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2533.4]
  assign _T_3232 = dat_rsp_p0_vld_w & dat_rsp_mask_w_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2537.4]
  assign _T_3233 = dat_rsp_p0_vld_w & dat_rsp_mask_w_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2541.4]
  assign _T_3234 = dat_rsp_p0_vld_w & dat_rsp_mask_w_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2545.4]
  assign _T_3235 = dat_rsp_p0_vld_w & dat_rsp_mask_w_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2549.4]
  assign _T_3236 = dat_rsp_p0_vld_w & dat_rsp_mask_w_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2553.4]
  assign _T_3237 = dat_rsp_p0_vld_w & dat_rsp_mask_w_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2557.4]
  assign _T_3238 = dat_rsp_p0_vld_w & dat_rsp_mask_w_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2561.4]
  assign _T_3239 = dat_rsp_p0_vld_w & dat_rsp_mask_w_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2565.4]
  assign _T_3240 = dat_rsp_p0_vld_w & dat_rsp_mask_w_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2569.4]
  assign _T_3241 = dat_rsp_p0_vld_w & dat_rsp_mask_w_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2573.4]
  assign _T_3242 = dat_rsp_p0_vld_w & dat_rsp_mask_w_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1168:34:@2577.4]
  assign _T_4044 = is_winograd_d1[20]; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:38:@2780.4]
  assign dat_out_data_0 = _T_4044 ? 8'h0 : dat_out_bypass_data_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_1 = _T_4044 ? 8'h0 : dat_out_bypass_data_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_2 = _T_4044 ? 8'h0 : dat_out_bypass_data_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_3 = _T_4044 ? 8'h0 : dat_out_bypass_data_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_4 = _T_4044 ? 8'h0 : dat_out_bypass_data_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_5 = _T_4044 ? 8'h0 : dat_out_bypass_data_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_6 = _T_4044 ? 8'h0 : dat_out_bypass_data_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_7 = _T_4044 ? 8'h0 : dat_out_bypass_data_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_8 = _T_4044 ? 8'h0 : dat_out_bypass_data_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_9 = _T_4044 ? 8'h0 : dat_out_bypass_data_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_10 = _T_4044 ? 8'h0 : dat_out_bypass_data_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_11 = _T_4044 ? 8'h0 : dat_out_bypass_data_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_12 = _T_4044 ? 8'h0 : dat_out_bypass_data_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_13 = _T_4044 ? 8'h0 : dat_out_bypass_data_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_14 = _T_4044 ? 8'h0 : dat_out_bypass_data_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_15 = _T_4044 ? 8'h0 : dat_out_bypass_data_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_16 = _T_4044 ? 8'h0 : dat_out_bypass_data_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_17 = _T_4044 ? 8'h0 : dat_out_bypass_data_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_18 = _T_4044 ? 8'h0 : dat_out_bypass_data_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_19 = _T_4044 ? 8'h0 : dat_out_bypass_data_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_20 = _T_4044 ? 8'h0 : dat_out_bypass_data_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_21 = _T_4044 ? 8'h0 : dat_out_bypass_data_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_22 = _T_4044 ? 8'h0 : dat_out_bypass_data_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_23 = _T_4044 ? 8'h0 : dat_out_bypass_data_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_24 = _T_4044 ? 8'h0 : dat_out_bypass_data_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_25 = _T_4044 ? 8'h0 : dat_out_bypass_data_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_26 = _T_4044 ? 8'h0 : dat_out_bypass_data_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_27 = _T_4044 ? 8'h0 : dat_out_bypass_data_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_28 = _T_4044 ? 8'h0 : dat_out_bypass_data_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_29 = _T_4044 ? 8'h0 : dat_out_bypass_data_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_30 = _T_4044 ? 8'h0 : dat_out_bypass_data_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_31 = _T_4044 ? 8'h0 : dat_out_bypass_data_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_32 = _T_4044 ? 8'h0 : dat_out_bypass_data_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_33 = _T_4044 ? 8'h0 : dat_out_bypass_data_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_34 = _T_4044 ? 8'h0 : dat_out_bypass_data_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_35 = _T_4044 ? 8'h0 : dat_out_bypass_data_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_36 = _T_4044 ? 8'h0 : dat_out_bypass_data_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_37 = _T_4044 ? 8'h0 : dat_out_bypass_data_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_38 = _T_4044 ? 8'h0 : dat_out_bypass_data_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_39 = _T_4044 ? 8'h0 : dat_out_bypass_data_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_40 = _T_4044 ? 8'h0 : dat_out_bypass_data_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_41 = _T_4044 ? 8'h0 : dat_out_bypass_data_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_42 = _T_4044 ? 8'h0 : dat_out_bypass_data_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_43 = _T_4044 ? 8'h0 : dat_out_bypass_data_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_44 = _T_4044 ? 8'h0 : dat_out_bypass_data_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_45 = _T_4044 ? 8'h0 : dat_out_bypass_data_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_46 = _T_4044 ? 8'h0 : dat_out_bypass_data_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_47 = _T_4044 ? 8'h0 : dat_out_bypass_data_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_48 = _T_4044 ? 8'h0 : dat_out_bypass_data_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_49 = _T_4044 ? 8'h0 : dat_out_bypass_data_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_50 = _T_4044 ? 8'h0 : dat_out_bypass_data_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_51 = _T_4044 ? 8'h0 : dat_out_bypass_data_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_52 = _T_4044 ? 8'h0 : dat_out_bypass_data_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_53 = _T_4044 ? 8'h0 : dat_out_bypass_data_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_54 = _T_4044 ? 8'h0 : dat_out_bypass_data_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_55 = _T_4044 ? 8'h0 : dat_out_bypass_data_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_56 = _T_4044 ? 8'h0 : dat_out_bypass_data_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_57 = _T_4044 ? 8'h0 : dat_out_bypass_data_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_58 = _T_4044 ? 8'h0 : dat_out_bypass_data_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_59 = _T_4044 ? 8'h0 : dat_out_bypass_data_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_60 = _T_4044 ? 8'h0 : dat_out_bypass_data_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_61 = _T_4044 ? 8'h0 : dat_out_bypass_data_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_62 = _T_4044 ? 8'h0 : dat_out_bypass_data_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign dat_out_data_63 = _T_4044 ? 8'h0 : dat_out_bypass_data_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1187:23:@2781.4]
  assign _T_4176 = ~ dat_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:24:@2782.4]
  assign _T_4311 = is_winograd_d1[21]; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:38:@2848.4]
  assign _T_4312_0 = _T_4311 ? 1'h0 : dat_out_bypass_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_1 = _T_4311 ? 1'h0 : dat_out_bypass_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_2 = _T_4311 ? 1'h0 : dat_out_bypass_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_3 = _T_4311 ? 1'h0 : dat_out_bypass_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_4 = _T_4311 ? 1'h0 : dat_out_bypass_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_5 = _T_4311 ? 1'h0 : dat_out_bypass_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_6 = _T_4311 ? 1'h0 : dat_out_bypass_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_7 = _T_4311 ? 1'h0 : dat_out_bypass_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_8 = _T_4311 ? 1'h0 : dat_out_bypass_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_9 = _T_4311 ? 1'h0 : dat_out_bypass_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_10 = _T_4311 ? 1'h0 : dat_out_bypass_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_11 = _T_4311 ? 1'h0 : dat_out_bypass_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_12 = _T_4311 ? 1'h0 : dat_out_bypass_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_13 = _T_4311 ? 1'h0 : dat_out_bypass_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_14 = _T_4311 ? 1'h0 : dat_out_bypass_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_15 = _T_4311 ? 1'h0 : dat_out_bypass_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_16 = _T_4311 ? 1'h0 : dat_out_bypass_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_17 = _T_4311 ? 1'h0 : dat_out_bypass_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_18 = _T_4311 ? 1'h0 : dat_out_bypass_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_19 = _T_4311 ? 1'h0 : dat_out_bypass_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_20 = _T_4311 ? 1'h0 : dat_out_bypass_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_21 = _T_4311 ? 1'h0 : dat_out_bypass_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_22 = _T_4311 ? 1'h0 : dat_out_bypass_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_23 = _T_4311 ? 1'h0 : dat_out_bypass_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_24 = _T_4311 ? 1'h0 : dat_out_bypass_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_25 = _T_4311 ? 1'h0 : dat_out_bypass_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_26 = _T_4311 ? 1'h0 : dat_out_bypass_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_27 = _T_4311 ? 1'h0 : dat_out_bypass_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_28 = _T_4311 ? 1'h0 : dat_out_bypass_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_29 = _T_4311 ? 1'h0 : dat_out_bypass_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_30 = _T_4311 ? 1'h0 : dat_out_bypass_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_31 = _T_4311 ? 1'h0 : dat_out_bypass_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_32 = _T_4311 ? 1'h0 : dat_out_bypass_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_33 = _T_4311 ? 1'h0 : dat_out_bypass_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_34 = _T_4311 ? 1'h0 : dat_out_bypass_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_35 = _T_4311 ? 1'h0 : dat_out_bypass_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_36 = _T_4311 ? 1'h0 : dat_out_bypass_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_37 = _T_4311 ? 1'h0 : dat_out_bypass_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_38 = _T_4311 ? 1'h0 : dat_out_bypass_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_39 = _T_4311 ? 1'h0 : dat_out_bypass_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_40 = _T_4311 ? 1'h0 : dat_out_bypass_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_41 = _T_4311 ? 1'h0 : dat_out_bypass_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_42 = _T_4311 ? 1'h0 : dat_out_bypass_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_43 = _T_4311 ? 1'h0 : dat_out_bypass_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_44 = _T_4311 ? 1'h0 : dat_out_bypass_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_45 = _T_4311 ? 1'h0 : dat_out_bypass_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_46 = _T_4311 ? 1'h0 : dat_out_bypass_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_47 = _T_4311 ? 1'h0 : dat_out_bypass_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_48 = _T_4311 ? 1'h0 : dat_out_bypass_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_49 = _T_4311 ? 1'h0 : dat_out_bypass_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_50 = _T_4311 ? 1'h0 : dat_out_bypass_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_51 = _T_4311 ? 1'h0 : dat_out_bypass_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_52 = _T_4311 ? 1'h0 : dat_out_bypass_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_53 = _T_4311 ? 1'h0 : dat_out_bypass_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_54 = _T_4311 ? 1'h0 : dat_out_bypass_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_55 = _T_4311 ? 1'h0 : dat_out_bypass_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_56 = _T_4311 ? 1'h0 : dat_out_bypass_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_57 = _T_4311 ? 1'h0 : dat_out_bypass_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_58 = _T_4311 ? 1'h0 : dat_out_bypass_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_59 = _T_4311 ? 1'h0 : dat_out_bypass_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_60 = _T_4311 ? 1'h0 : dat_out_bypass_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_61 = _T_4311 ? 1'h0 : dat_out_bypass_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_62 = _T_4311 ? 1'h0 : dat_out_bypass_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign _T_4312_63 = _T_4311 ? 1'h0 : dat_out_bypass_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1189:23:@2849.4]
  assign dat_out_mask_0 = _T_4176 ? 1'h0 : _T_4312_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_1 = _T_4176 ? 1'h0 : _T_4312_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_2 = _T_4176 ? 1'h0 : _T_4312_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_3 = _T_4176 ? 1'h0 : _T_4312_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_4 = _T_4176 ? 1'h0 : _T_4312_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_5 = _T_4176 ? 1'h0 : _T_4312_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_6 = _T_4176 ? 1'h0 : _T_4312_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_7 = _T_4176 ? 1'h0 : _T_4312_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_8 = _T_4176 ? 1'h0 : _T_4312_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_9 = _T_4176 ? 1'h0 : _T_4312_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_10 = _T_4176 ? 1'h0 : _T_4312_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_11 = _T_4176 ? 1'h0 : _T_4312_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_12 = _T_4176 ? 1'h0 : _T_4312_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_13 = _T_4176 ? 1'h0 : _T_4312_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_14 = _T_4176 ? 1'h0 : _T_4312_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_15 = _T_4176 ? 1'h0 : _T_4312_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_16 = _T_4176 ? 1'h0 : _T_4312_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_17 = _T_4176 ? 1'h0 : _T_4312_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_18 = _T_4176 ? 1'h0 : _T_4312_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_19 = _T_4176 ? 1'h0 : _T_4312_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_20 = _T_4176 ? 1'h0 : _T_4312_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_21 = _T_4176 ? 1'h0 : _T_4312_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_22 = _T_4176 ? 1'h0 : _T_4312_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_23 = _T_4176 ? 1'h0 : _T_4312_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_24 = _T_4176 ? 1'h0 : _T_4312_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_25 = _T_4176 ? 1'h0 : _T_4312_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_26 = _T_4176 ? 1'h0 : _T_4312_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_27 = _T_4176 ? 1'h0 : _T_4312_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_28 = _T_4176 ? 1'h0 : _T_4312_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_29 = _T_4176 ? 1'h0 : _T_4312_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_30 = _T_4176 ? 1'h0 : _T_4312_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_31 = _T_4176 ? 1'h0 : _T_4312_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_32 = _T_4176 ? 1'h0 : _T_4312_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_33 = _T_4176 ? 1'h0 : _T_4312_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_34 = _T_4176 ? 1'h0 : _T_4312_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_35 = _T_4176 ? 1'h0 : _T_4312_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_36 = _T_4176 ? 1'h0 : _T_4312_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_37 = _T_4176 ? 1'h0 : _T_4312_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_38 = _T_4176 ? 1'h0 : _T_4312_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_39 = _T_4176 ? 1'h0 : _T_4312_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_40 = _T_4176 ? 1'h0 : _T_4312_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_41 = _T_4176 ? 1'h0 : _T_4312_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_42 = _T_4176 ? 1'h0 : _T_4312_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_43 = _T_4176 ? 1'h0 : _T_4312_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_44 = _T_4176 ? 1'h0 : _T_4312_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_45 = _T_4176 ? 1'h0 : _T_4312_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_46 = _T_4176 ? 1'h0 : _T_4312_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_47 = _T_4176 ? 1'h0 : _T_4312_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_48 = _T_4176 ? 1'h0 : _T_4312_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_49 = _T_4176 ? 1'h0 : _T_4312_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_50 = _T_4176 ? 1'h0 : _T_4312_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_51 = _T_4176 ? 1'h0 : _T_4312_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_52 = _T_4176 ? 1'h0 : _T_4312_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_53 = _T_4176 ? 1'h0 : _T_4312_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_54 = _T_4176 ? 1'h0 : _T_4312_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_55 = _T_4176 ? 1'h0 : _T_4312_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_56 = _T_4176 ? 1'h0 : _T_4312_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_57 = _T_4176 ? 1'h0 : _T_4312_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_58 = _T_4176 ? 1'h0 : _T_4312_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_59 = _T_4176 ? 1'h0 : _T_4312_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_60 = _T_4176 ? 1'h0 : _T_4312_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_61 = _T_4176 ? 1'h0 : _T_4312_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_62 = _T_4176 ? 1'h0 : _T_4312_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign dat_out_mask_63 = _T_4176 ? 1'h0 : _T_4312_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1188:23:@2850.4]
  assign _T_4575 = dat_out_pvld | dl_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:19:@2852.4]
  assign _GEN_294 = _T_4575 ? dat_out_mask_0 : dl_out_mask_0; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_295 = _T_4575 ? dat_out_mask_1 : dl_out_mask_1; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_296 = _T_4575 ? dat_out_mask_2 : dl_out_mask_2; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_297 = _T_4575 ? dat_out_mask_3 : dl_out_mask_3; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_298 = _T_4575 ? dat_out_mask_4 : dl_out_mask_4; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_299 = _T_4575 ? dat_out_mask_5 : dl_out_mask_5; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_300 = _T_4575 ? dat_out_mask_6 : dl_out_mask_6; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_301 = _T_4575 ? dat_out_mask_7 : dl_out_mask_7; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_302 = _T_4575 ? dat_out_mask_8 : dl_out_mask_8; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_303 = _T_4575 ? dat_out_mask_9 : dl_out_mask_9; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_304 = _T_4575 ? dat_out_mask_10 : dl_out_mask_10; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_305 = _T_4575 ? dat_out_mask_11 : dl_out_mask_11; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_306 = _T_4575 ? dat_out_mask_12 : dl_out_mask_12; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_307 = _T_4575 ? dat_out_mask_13 : dl_out_mask_13; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_308 = _T_4575 ? dat_out_mask_14 : dl_out_mask_14; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_309 = _T_4575 ? dat_out_mask_15 : dl_out_mask_15; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_310 = _T_4575 ? dat_out_mask_16 : dl_out_mask_16; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_311 = _T_4575 ? dat_out_mask_17 : dl_out_mask_17; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_312 = _T_4575 ? dat_out_mask_18 : dl_out_mask_18; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_313 = _T_4575 ? dat_out_mask_19 : dl_out_mask_19; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_314 = _T_4575 ? dat_out_mask_20 : dl_out_mask_20; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_315 = _T_4575 ? dat_out_mask_21 : dl_out_mask_21; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_316 = _T_4575 ? dat_out_mask_22 : dl_out_mask_22; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_317 = _T_4575 ? dat_out_mask_23 : dl_out_mask_23; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_318 = _T_4575 ? dat_out_mask_24 : dl_out_mask_24; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_319 = _T_4575 ? dat_out_mask_25 : dl_out_mask_25; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_320 = _T_4575 ? dat_out_mask_26 : dl_out_mask_26; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_321 = _T_4575 ? dat_out_mask_27 : dl_out_mask_27; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_322 = _T_4575 ? dat_out_mask_28 : dl_out_mask_28; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_323 = _T_4575 ? dat_out_mask_29 : dl_out_mask_29; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_324 = _T_4575 ? dat_out_mask_30 : dl_out_mask_30; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_325 = _T_4575 ? dat_out_mask_31 : dl_out_mask_31; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_326 = _T_4575 ? dat_out_mask_32 : dl_out_mask_32; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_327 = _T_4575 ? dat_out_mask_33 : dl_out_mask_33; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_328 = _T_4575 ? dat_out_mask_34 : dl_out_mask_34; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_329 = _T_4575 ? dat_out_mask_35 : dl_out_mask_35; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_330 = _T_4575 ? dat_out_mask_36 : dl_out_mask_36; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_331 = _T_4575 ? dat_out_mask_37 : dl_out_mask_37; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_332 = _T_4575 ? dat_out_mask_38 : dl_out_mask_38; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_333 = _T_4575 ? dat_out_mask_39 : dl_out_mask_39; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_334 = _T_4575 ? dat_out_mask_40 : dl_out_mask_40; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_335 = _T_4575 ? dat_out_mask_41 : dl_out_mask_41; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_336 = _T_4575 ? dat_out_mask_42 : dl_out_mask_42; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_337 = _T_4575 ? dat_out_mask_43 : dl_out_mask_43; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_338 = _T_4575 ? dat_out_mask_44 : dl_out_mask_44; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_339 = _T_4575 ? dat_out_mask_45 : dl_out_mask_45; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_340 = _T_4575 ? dat_out_mask_46 : dl_out_mask_46; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_341 = _T_4575 ? dat_out_mask_47 : dl_out_mask_47; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_342 = _T_4575 ? dat_out_mask_48 : dl_out_mask_48; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_343 = _T_4575 ? dat_out_mask_49 : dl_out_mask_49; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_344 = _T_4575 ? dat_out_mask_50 : dl_out_mask_50; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_345 = _T_4575 ? dat_out_mask_51 : dl_out_mask_51; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_346 = _T_4575 ? dat_out_mask_52 : dl_out_mask_52; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_347 = _T_4575 ? dat_out_mask_53 : dl_out_mask_53; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_348 = _T_4575 ? dat_out_mask_54 : dl_out_mask_54; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_349 = _T_4575 ? dat_out_mask_55 : dl_out_mask_55; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_350 = _T_4575 ? dat_out_mask_56 : dl_out_mask_56; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_351 = _T_4575 ? dat_out_mask_57 : dl_out_mask_57; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_352 = _T_4575 ? dat_out_mask_58 : dl_out_mask_58; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_353 = _T_4575 ? dat_out_mask_59 : dl_out_mask_59; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_354 = _T_4575 ? dat_out_mask_60 : dl_out_mask_60; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_355 = _T_4575 ? dat_out_mask_61 : dl_out_mask_61; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_356 = _T_4575 ? dat_out_mask_62 : dl_out_mask_62; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_357 = _T_4575 ? dat_out_mask_63 : dl_out_mask_63; // @[NV_NVDLA_CSC_dl_for_check.scala 1192:33:@2853.4]
  assign _GEN_358 = dat_out_pvld ? dat_out_flag : dl_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1195:19:@2919.4]
  assign _T_4578 = ~ dl_out_pvld; // @[NV_NVDLA_CSC_dl_for_check.scala 1209:27:@3116.4]
  assign sc2mac_dat_pd_w = _T_4578 ? 9'h0 : dl_out_flag; // @[NV_NVDLA_CSC_dl_for_check.scala 1209:26:@3117.4]
  assign _T_4587 = dl_out_pvld | dl_out_pvld_d1; // @[NV_NVDLA_CSC_dl_for_check.scala 1213:80:@3124.4]
  assign _GEN_423 = _T_4587 ? sc2mac_dat_pd_w : _T_4589; // @[Reg.scala 20:19:@3126.4]
  assign _GEN_424 = _T_4587 ? sc2mac_dat_pd_w : _T_4593; // @[Reg.scala 20:19:@3132.4]
  assign _GEN_425 = _T_4587 ? dl_out_mask_0 : _T_4861_0; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_426 = _T_4587 ? dl_out_mask_1 : _T_4861_1; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_427 = _T_4587 ? dl_out_mask_2 : _T_4861_2; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_428 = _T_4587 ? dl_out_mask_3 : _T_4861_3; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_429 = _T_4587 ? dl_out_mask_4 : _T_4861_4; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_430 = _T_4587 ? dl_out_mask_5 : _T_4861_5; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_431 = _T_4587 ? dl_out_mask_6 : _T_4861_6; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_432 = _T_4587 ? dl_out_mask_7 : _T_4861_7; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_433 = _T_4587 ? dl_out_mask_8 : _T_4861_8; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_434 = _T_4587 ? dl_out_mask_9 : _T_4861_9; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_435 = _T_4587 ? dl_out_mask_10 : _T_4861_10; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_436 = _T_4587 ? dl_out_mask_11 : _T_4861_11; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_437 = _T_4587 ? dl_out_mask_12 : _T_4861_12; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_438 = _T_4587 ? dl_out_mask_13 : _T_4861_13; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_439 = _T_4587 ? dl_out_mask_14 : _T_4861_14; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_440 = _T_4587 ? dl_out_mask_15 : _T_4861_15; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_441 = _T_4587 ? dl_out_mask_16 : _T_4861_16; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_442 = _T_4587 ? dl_out_mask_17 : _T_4861_17; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_443 = _T_4587 ? dl_out_mask_18 : _T_4861_18; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_444 = _T_4587 ? dl_out_mask_19 : _T_4861_19; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_445 = _T_4587 ? dl_out_mask_20 : _T_4861_20; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_446 = _T_4587 ? dl_out_mask_21 : _T_4861_21; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_447 = _T_4587 ? dl_out_mask_22 : _T_4861_22; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_448 = _T_4587 ? dl_out_mask_23 : _T_4861_23; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_449 = _T_4587 ? dl_out_mask_24 : _T_4861_24; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_450 = _T_4587 ? dl_out_mask_25 : _T_4861_25; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_451 = _T_4587 ? dl_out_mask_26 : _T_4861_26; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_452 = _T_4587 ? dl_out_mask_27 : _T_4861_27; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_453 = _T_4587 ? dl_out_mask_28 : _T_4861_28; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_454 = _T_4587 ? dl_out_mask_29 : _T_4861_29; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_455 = _T_4587 ? dl_out_mask_30 : _T_4861_30; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_456 = _T_4587 ? dl_out_mask_31 : _T_4861_31; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_457 = _T_4587 ? dl_out_mask_32 : _T_4861_32; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_458 = _T_4587 ? dl_out_mask_33 : _T_4861_33; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_459 = _T_4587 ? dl_out_mask_34 : _T_4861_34; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_460 = _T_4587 ? dl_out_mask_35 : _T_4861_35; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_461 = _T_4587 ? dl_out_mask_36 : _T_4861_36; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_462 = _T_4587 ? dl_out_mask_37 : _T_4861_37; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_463 = _T_4587 ? dl_out_mask_38 : _T_4861_38; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_464 = _T_4587 ? dl_out_mask_39 : _T_4861_39; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_465 = _T_4587 ? dl_out_mask_40 : _T_4861_40; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_466 = _T_4587 ? dl_out_mask_41 : _T_4861_41; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_467 = _T_4587 ? dl_out_mask_42 : _T_4861_42; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_468 = _T_4587 ? dl_out_mask_43 : _T_4861_43; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_469 = _T_4587 ? dl_out_mask_44 : _T_4861_44; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_470 = _T_4587 ? dl_out_mask_45 : _T_4861_45; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_471 = _T_4587 ? dl_out_mask_46 : _T_4861_46; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_472 = _T_4587 ? dl_out_mask_47 : _T_4861_47; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_473 = _T_4587 ? dl_out_mask_48 : _T_4861_48; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_474 = _T_4587 ? dl_out_mask_49 : _T_4861_49; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_475 = _T_4587 ? dl_out_mask_50 : _T_4861_50; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_476 = _T_4587 ? dl_out_mask_51 : _T_4861_51; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_477 = _T_4587 ? dl_out_mask_52 : _T_4861_52; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_478 = _T_4587 ? dl_out_mask_53 : _T_4861_53; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_479 = _T_4587 ? dl_out_mask_54 : _T_4861_54; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_480 = _T_4587 ? dl_out_mask_55 : _T_4861_55; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_481 = _T_4587 ? dl_out_mask_56 : _T_4861_56; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_482 = _T_4587 ? dl_out_mask_57 : _T_4861_57; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_483 = _T_4587 ? dl_out_mask_58 : _T_4861_58; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_484 = _T_4587 ? dl_out_mask_59 : _T_4861_59; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_485 = _T_4587 ? dl_out_mask_60 : _T_4861_60; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_486 = _T_4587 ? dl_out_mask_61 : _T_4861_61; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_487 = _T_4587 ? dl_out_mask_62 : _T_4861_62; // @[Reg.scala 20:19:@3203.4]
  assign _GEN_488 = _T_4587 ? dl_out_mask_63 : _T_4861_63; // @[Reg.scala 20:19:@3203.4]
  assign _T_5064 = {_T_4861_7,_T_4861_6,_T_4861_5,_T_4861_4,_T_4861_3,_T_4861_2,_T_4861_1,_T_4861_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3275.4]
  assign _T_5072 = {_T_4861_15,_T_4861_14,_T_4861_13,_T_4861_12,_T_4861_11,_T_4861_10,_T_4861_9,_T_4861_8,_T_5064}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3283.4]
  assign _T_5079 = {_T_4861_23,_T_4861_22,_T_4861_21,_T_4861_20,_T_4861_19,_T_4861_18,_T_4861_17,_T_4861_16}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3290.4]
  assign _T_5088 = {_T_4861_31,_T_4861_30,_T_4861_29,_T_4861_28,_T_4861_27,_T_4861_26,_T_4861_25,_T_4861_24,_T_5079,_T_5072}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3299.4]
  assign _T_5095 = {_T_4861_39,_T_4861_38,_T_4861_37,_T_4861_36,_T_4861_35,_T_4861_34,_T_4861_33,_T_4861_32}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3306.4]
  assign _T_5103 = {_T_4861_47,_T_4861_46,_T_4861_45,_T_4861_44,_T_4861_43,_T_4861_42,_T_4861_41,_T_4861_40,_T_5095}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3314.4]
  assign _T_5110 = {_T_4861_55,_T_4861_54,_T_4861_53,_T_4861_52,_T_4861_51,_T_4861_50,_T_4861_49,_T_4861_48}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3321.4]
  assign _T_5119 = {_T_4861_63,_T_4861_62,_T_4861_61,_T_4861_60,_T_4861_59,_T_4861_58,_T_4861_57,_T_4861_56,_T_5110,_T_5103}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:122:@3330.4]
  assign _GEN_489 = _T_4587 ? dl_out_mask_0 : _T_5388_0; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_490 = _T_4587 ? dl_out_mask_1 : _T_5388_1; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_491 = _T_4587 ? dl_out_mask_2 : _T_5388_2; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_492 = _T_4587 ? dl_out_mask_3 : _T_5388_3; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_493 = _T_4587 ? dl_out_mask_4 : _T_5388_4; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_494 = _T_4587 ? dl_out_mask_5 : _T_5388_5; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_495 = _T_4587 ? dl_out_mask_6 : _T_5388_6; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_496 = _T_4587 ? dl_out_mask_7 : _T_5388_7; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_497 = _T_4587 ? dl_out_mask_8 : _T_5388_8; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_498 = _T_4587 ? dl_out_mask_9 : _T_5388_9; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_499 = _T_4587 ? dl_out_mask_10 : _T_5388_10; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_500 = _T_4587 ? dl_out_mask_11 : _T_5388_11; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_501 = _T_4587 ? dl_out_mask_12 : _T_5388_12; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_502 = _T_4587 ? dl_out_mask_13 : _T_5388_13; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_503 = _T_4587 ? dl_out_mask_14 : _T_5388_14; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_504 = _T_4587 ? dl_out_mask_15 : _T_5388_15; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_505 = _T_4587 ? dl_out_mask_16 : _T_5388_16; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_506 = _T_4587 ? dl_out_mask_17 : _T_5388_17; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_507 = _T_4587 ? dl_out_mask_18 : _T_5388_18; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_508 = _T_4587 ? dl_out_mask_19 : _T_5388_19; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_509 = _T_4587 ? dl_out_mask_20 : _T_5388_20; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_510 = _T_4587 ? dl_out_mask_21 : _T_5388_21; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_511 = _T_4587 ? dl_out_mask_22 : _T_5388_22; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_512 = _T_4587 ? dl_out_mask_23 : _T_5388_23; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_513 = _T_4587 ? dl_out_mask_24 : _T_5388_24; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_514 = _T_4587 ? dl_out_mask_25 : _T_5388_25; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_515 = _T_4587 ? dl_out_mask_26 : _T_5388_26; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_516 = _T_4587 ? dl_out_mask_27 : _T_5388_27; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_517 = _T_4587 ? dl_out_mask_28 : _T_5388_28; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_518 = _T_4587 ? dl_out_mask_29 : _T_5388_29; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_519 = _T_4587 ? dl_out_mask_30 : _T_5388_30; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_520 = _T_4587 ? dl_out_mask_31 : _T_5388_31; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_521 = _T_4587 ? dl_out_mask_32 : _T_5388_32; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_522 = _T_4587 ? dl_out_mask_33 : _T_5388_33; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_523 = _T_4587 ? dl_out_mask_34 : _T_5388_34; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_524 = _T_4587 ? dl_out_mask_35 : _T_5388_35; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_525 = _T_4587 ? dl_out_mask_36 : _T_5388_36; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_526 = _T_4587 ? dl_out_mask_37 : _T_5388_37; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_527 = _T_4587 ? dl_out_mask_38 : _T_5388_38; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_528 = _T_4587 ? dl_out_mask_39 : _T_5388_39; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_529 = _T_4587 ? dl_out_mask_40 : _T_5388_40; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_530 = _T_4587 ? dl_out_mask_41 : _T_5388_41; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_531 = _T_4587 ? dl_out_mask_42 : _T_5388_42; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_532 = _T_4587 ? dl_out_mask_43 : _T_5388_43; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_533 = _T_4587 ? dl_out_mask_44 : _T_5388_44; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_534 = _T_4587 ? dl_out_mask_45 : _T_5388_45; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_535 = _T_4587 ? dl_out_mask_46 : _T_5388_46; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_536 = _T_4587 ? dl_out_mask_47 : _T_5388_47; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_537 = _T_4587 ? dl_out_mask_48 : _T_5388_48; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_538 = _T_4587 ? dl_out_mask_49 : _T_5388_49; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_539 = _T_4587 ? dl_out_mask_50 : _T_5388_50; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_540 = _T_4587 ? dl_out_mask_51 : _T_5388_51; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_541 = _T_4587 ? dl_out_mask_52 : _T_5388_52; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_542 = _T_4587 ? dl_out_mask_53 : _T_5388_53; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_543 = _T_4587 ? dl_out_mask_54 : _T_5388_54; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_544 = _T_4587 ? dl_out_mask_55 : _T_5388_55; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_545 = _T_4587 ? dl_out_mask_56 : _T_5388_56; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_546 = _T_4587 ? dl_out_mask_57 : _T_5388_57; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_547 = _T_4587 ? dl_out_mask_58 : _T_5388_58; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_548 = _T_4587 ? dl_out_mask_59 : _T_5388_59; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_549 = _T_4587 ? dl_out_mask_60 : _T_5388_60; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_550 = _T_4587 ? dl_out_mask_61 : _T_5388_61; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_551 = _T_4587 ? dl_out_mask_62 : _T_5388_62; // @[Reg.scala 20:19:@3400.4]
  assign _GEN_552 = _T_4587 ? dl_out_mask_63 : _T_5388_63; // @[Reg.scala 20:19:@3400.4]
  assign _T_5591 = {_T_5388_7,_T_5388_6,_T_5388_5,_T_5388_4,_T_5388_3,_T_5388_2,_T_5388_1,_T_5388_0}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3472.4]
  assign _T_5599 = {_T_5388_15,_T_5388_14,_T_5388_13,_T_5388_12,_T_5388_11,_T_5388_10,_T_5388_9,_T_5388_8,_T_5591}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3480.4]
  assign _T_5606 = {_T_5388_23,_T_5388_22,_T_5388_21,_T_5388_20,_T_5388_19,_T_5388_18,_T_5388_17,_T_5388_16}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3487.4]
  assign _T_5615 = {_T_5388_31,_T_5388_30,_T_5388_29,_T_5388_28,_T_5388_27,_T_5388_26,_T_5388_25,_T_5388_24,_T_5606,_T_5599}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3496.4]
  assign _T_5622 = {_T_5388_39,_T_5388_38,_T_5388_37,_T_5388_36,_T_5388_35,_T_5388_34,_T_5388_33,_T_5388_32}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3503.4]
  assign _T_5630 = {_T_5388_47,_T_5388_46,_T_5388_45,_T_5388_44,_T_5388_43,_T_5388_42,_T_5388_41,_T_5388_40,_T_5622}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3511.4]
  assign _T_5637 = {_T_5388_55,_T_5388_54,_T_5388_53,_T_5388_52,_T_5388_51,_T_5388_50,_T_5388_49,_T_5388_48}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3518.4]
  assign _T_5646 = {_T_5388_63,_T_5388_62,_T_5388_61,_T_5388_60,_T_5388_59,_T_5388_58,_T_5388_57,_T_5388_56,_T_5637,_T_5630}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:122:@3527.4]
  assign io_sc2cdma_dat_updt_valid = _T_653; // @[NV_NVDLA_CSC_dl_for_check.scala 319:27:@340.4]
  assign io_sc2cdma_dat_updt_bits_entries = _T_659; // @[NV_NVDLA_CSC_dl_for_check.scala 321:34:@350.4]
  assign io_sc2cdma_dat_updt_bits_slices = _T_656; // @[NV_NVDLA_CSC_dl_for_check.scala 320:33:@345.4]
  assign io_sc2buf_dat_rd_addr_valid = sc2buf_dat_rd_en_out; // @[NV_NVDLA_CSC_dl_for_check.scala 742:29:@951.4]
  assign io_sc2buf_dat_rd_addr_bits = sc2buf_dat_rd_addr_out[12:0]; // @[NV_NVDLA_CSC_dl_for_check.scala 743:28:@952.4]
  assign io_sc2mac_dat_a_pvld = _T_4582; // @[NV_NVDLA_CSC_dl_for_check.scala 1211:22:@3120.4]
  assign io_sc2mac_dat_a_mask = {_T_5119,_T_5088}; // @[NV_NVDLA_CSC_dl_for_check.scala 1215:22:@3332.4]
  assign io_sc2mac_dat_a_data_0 = _T_5649; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3534.4]
  assign io_sc2mac_dat_a_data_1 = _T_5653; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3544.4]
  assign io_sc2mac_dat_a_data_2 = _T_5657; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3554.4]
  assign io_sc2mac_dat_a_data_3 = _T_5661; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3564.4]
  assign io_sc2mac_dat_a_data_4 = _T_5665; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3574.4]
  assign io_sc2mac_dat_a_data_5 = _T_5669; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3584.4]
  assign io_sc2mac_dat_a_data_6 = _T_5673; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3594.4]
  assign io_sc2mac_dat_a_data_7 = _T_5677; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3604.4]
  assign io_sc2mac_dat_a_data_8 = _T_5681; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3614.4]
  assign io_sc2mac_dat_a_data_9 = _T_5685; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3624.4]
  assign io_sc2mac_dat_a_data_10 = _T_5689; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3634.4]
  assign io_sc2mac_dat_a_data_11 = _T_5693; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3644.4]
  assign io_sc2mac_dat_a_data_12 = _T_5697; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3654.4]
  assign io_sc2mac_dat_a_data_13 = _T_5701; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3664.4]
  assign io_sc2mac_dat_a_data_14 = _T_5705; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3674.4]
  assign io_sc2mac_dat_a_data_15 = _T_5709; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3684.4]
  assign io_sc2mac_dat_a_data_16 = _T_5713; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3694.4]
  assign io_sc2mac_dat_a_data_17 = _T_5717; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3704.4]
  assign io_sc2mac_dat_a_data_18 = _T_5721; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3714.4]
  assign io_sc2mac_dat_a_data_19 = _T_5725; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3724.4]
  assign io_sc2mac_dat_a_data_20 = _T_5729; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3734.4]
  assign io_sc2mac_dat_a_data_21 = _T_5733; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3744.4]
  assign io_sc2mac_dat_a_data_22 = _T_5737; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3754.4]
  assign io_sc2mac_dat_a_data_23 = _T_5741; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3764.4]
  assign io_sc2mac_dat_a_data_24 = _T_5745; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3774.4]
  assign io_sc2mac_dat_a_data_25 = _T_5749; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3784.4]
  assign io_sc2mac_dat_a_data_26 = _T_5753; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3794.4]
  assign io_sc2mac_dat_a_data_27 = _T_5757; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3804.4]
  assign io_sc2mac_dat_a_data_28 = _T_5761; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3814.4]
  assign io_sc2mac_dat_a_data_29 = _T_5765; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3824.4]
  assign io_sc2mac_dat_a_data_30 = _T_5769; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3834.4]
  assign io_sc2mac_dat_a_data_31 = _T_5773; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3844.4]
  assign io_sc2mac_dat_a_data_32 = _T_5777; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3854.4]
  assign io_sc2mac_dat_a_data_33 = _T_5781; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3864.4]
  assign io_sc2mac_dat_a_data_34 = _T_5785; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3874.4]
  assign io_sc2mac_dat_a_data_35 = _T_5789; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3884.4]
  assign io_sc2mac_dat_a_data_36 = _T_5793; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3894.4]
  assign io_sc2mac_dat_a_data_37 = _T_5797; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3904.4]
  assign io_sc2mac_dat_a_data_38 = _T_5801; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3914.4]
  assign io_sc2mac_dat_a_data_39 = _T_5805; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3924.4]
  assign io_sc2mac_dat_a_data_40 = _T_5809; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3934.4]
  assign io_sc2mac_dat_a_data_41 = _T_5813; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3944.4]
  assign io_sc2mac_dat_a_data_42 = _T_5817; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3954.4]
  assign io_sc2mac_dat_a_data_43 = _T_5821; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3964.4]
  assign io_sc2mac_dat_a_data_44 = _T_5825; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3974.4]
  assign io_sc2mac_dat_a_data_45 = _T_5829; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3984.4]
  assign io_sc2mac_dat_a_data_46 = _T_5833; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@3994.4]
  assign io_sc2mac_dat_a_data_47 = _T_5837; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4004.4]
  assign io_sc2mac_dat_a_data_48 = _T_5841; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4014.4]
  assign io_sc2mac_dat_a_data_49 = _T_5845; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4024.4]
  assign io_sc2mac_dat_a_data_50 = _T_5849; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4034.4]
  assign io_sc2mac_dat_a_data_51 = _T_5853; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4044.4]
  assign io_sc2mac_dat_a_data_52 = _T_5857; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4054.4]
  assign io_sc2mac_dat_a_data_53 = _T_5861; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4064.4]
  assign io_sc2mac_dat_a_data_54 = _T_5865; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4074.4]
  assign io_sc2mac_dat_a_data_55 = _T_5869; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4084.4]
  assign io_sc2mac_dat_a_data_56 = _T_5873; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4094.4]
  assign io_sc2mac_dat_a_data_57 = _T_5877; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4104.4]
  assign io_sc2mac_dat_a_data_58 = _T_5881; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4114.4]
  assign io_sc2mac_dat_a_data_59 = _T_5885; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4124.4]
  assign io_sc2mac_dat_a_data_60 = _T_5889; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4134.4]
  assign io_sc2mac_dat_a_data_61 = _T_5893; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4144.4]
  assign io_sc2mac_dat_a_data_62 = _T_5897; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4154.4]
  assign io_sc2mac_dat_a_data_63 = _T_5901; // @[NV_NVDLA_CSC_dl_for_check.scala 1218:29:@4164.4]
  assign io_sc2mac_dat_a_pd = _T_4589; // @[NV_NVDLA_CSC_dl_for_check.scala 1213:20:@3129.4]
  assign io_sc2mac_dat_b_pvld = _T_4585; // @[NV_NVDLA_CSC_dl_for_check.scala 1212:22:@3123.4]
  assign io_sc2mac_dat_b_mask = {_T_5646,_T_5615}; // @[NV_NVDLA_CSC_dl_for_check.scala 1216:22:@3529.4]
  assign io_sc2mac_dat_b_data_0 = _T_5651; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3539.4]
  assign io_sc2mac_dat_b_data_1 = _T_5655; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3549.4]
  assign io_sc2mac_dat_b_data_2 = _T_5659; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3559.4]
  assign io_sc2mac_dat_b_data_3 = _T_5663; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3569.4]
  assign io_sc2mac_dat_b_data_4 = _T_5667; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3579.4]
  assign io_sc2mac_dat_b_data_5 = _T_5671; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3589.4]
  assign io_sc2mac_dat_b_data_6 = _T_5675; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3599.4]
  assign io_sc2mac_dat_b_data_7 = _T_5679; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3609.4]
  assign io_sc2mac_dat_b_data_8 = _T_5683; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3619.4]
  assign io_sc2mac_dat_b_data_9 = _T_5687; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3629.4]
  assign io_sc2mac_dat_b_data_10 = _T_5691; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3639.4]
  assign io_sc2mac_dat_b_data_11 = _T_5695; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3649.4]
  assign io_sc2mac_dat_b_data_12 = _T_5699; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3659.4]
  assign io_sc2mac_dat_b_data_13 = _T_5703; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3669.4]
  assign io_sc2mac_dat_b_data_14 = _T_5707; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3679.4]
  assign io_sc2mac_dat_b_data_15 = _T_5711; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3689.4]
  assign io_sc2mac_dat_b_data_16 = _T_5715; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3699.4]
  assign io_sc2mac_dat_b_data_17 = _T_5719; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3709.4]
  assign io_sc2mac_dat_b_data_18 = _T_5723; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3719.4]
  assign io_sc2mac_dat_b_data_19 = _T_5727; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3729.4]
  assign io_sc2mac_dat_b_data_20 = _T_5731; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3739.4]
  assign io_sc2mac_dat_b_data_21 = _T_5735; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3749.4]
  assign io_sc2mac_dat_b_data_22 = _T_5739; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3759.4]
  assign io_sc2mac_dat_b_data_23 = _T_5743; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3769.4]
  assign io_sc2mac_dat_b_data_24 = _T_5747; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3779.4]
  assign io_sc2mac_dat_b_data_25 = _T_5751; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3789.4]
  assign io_sc2mac_dat_b_data_26 = _T_5755; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3799.4]
  assign io_sc2mac_dat_b_data_27 = _T_5759; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3809.4]
  assign io_sc2mac_dat_b_data_28 = _T_5763; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3819.4]
  assign io_sc2mac_dat_b_data_29 = _T_5767; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3829.4]
  assign io_sc2mac_dat_b_data_30 = _T_5771; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3839.4]
  assign io_sc2mac_dat_b_data_31 = _T_5775; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3849.4]
  assign io_sc2mac_dat_b_data_32 = _T_5779; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3859.4]
  assign io_sc2mac_dat_b_data_33 = _T_5783; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3869.4]
  assign io_sc2mac_dat_b_data_34 = _T_5787; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3879.4]
  assign io_sc2mac_dat_b_data_35 = _T_5791; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3889.4]
  assign io_sc2mac_dat_b_data_36 = _T_5795; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3899.4]
  assign io_sc2mac_dat_b_data_37 = _T_5799; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3909.4]
  assign io_sc2mac_dat_b_data_38 = _T_5803; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3919.4]
  assign io_sc2mac_dat_b_data_39 = _T_5807; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3929.4]
  assign io_sc2mac_dat_b_data_40 = _T_5811; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3939.4]
  assign io_sc2mac_dat_b_data_41 = _T_5815; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3949.4]
  assign io_sc2mac_dat_b_data_42 = _T_5819; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3959.4]
  assign io_sc2mac_dat_b_data_43 = _T_5823; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3969.4]
  assign io_sc2mac_dat_b_data_44 = _T_5827; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3979.4]
  assign io_sc2mac_dat_b_data_45 = _T_5831; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3989.4]
  assign io_sc2mac_dat_b_data_46 = _T_5835; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@3999.4]
  assign io_sc2mac_dat_b_data_47 = _T_5839; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4009.4]
  assign io_sc2mac_dat_b_data_48 = _T_5843; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4019.4]
  assign io_sc2mac_dat_b_data_49 = _T_5847; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4029.4]
  assign io_sc2mac_dat_b_data_50 = _T_5851; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4039.4]
  assign io_sc2mac_dat_b_data_51 = _T_5855; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4049.4]
  assign io_sc2mac_dat_b_data_52 = _T_5859; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4059.4]
  assign io_sc2mac_dat_b_data_53 = _T_5863; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4069.4]
  assign io_sc2mac_dat_b_data_54 = _T_5867; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4079.4]
  assign io_sc2mac_dat_b_data_55 = _T_5871; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4089.4]
  assign io_sc2mac_dat_b_data_56 = _T_5875; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4099.4]
  assign io_sc2mac_dat_b_data_57 = _T_5879; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4109.4]
  assign io_sc2mac_dat_b_data_58 = _T_5883; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4119.4]
  assign io_sc2mac_dat_b_data_59 = _T_5887; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4129.4]
  assign io_sc2mac_dat_b_data_60 = _T_5891; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4139.4]
  assign io_sc2mac_dat_b_data_61 = _T_5895; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4149.4]
  assign io_sc2mac_dat_b_data_62 = _T_5899; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4159.4]
  assign io_sc2mac_dat_b_data_63 = _T_5903; // @[NV_NVDLA_CSC_dl_for_check.scala 1219:29:@4169.4]
  assign io_sc2mac_dat_b_pd = _T_4593; // @[NV_NVDLA_CSC_dl_for_check.scala 1214:20:@3135.4]
  assign io_slcg_wg_en = 1'h0; // @[NV_NVDLA_CSC_dl_for_check.scala 260:15:@261.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  layer_st_d1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  data_batch = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  rls_slices = _RAND_2[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  h_offset_slice = _RAND_3[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  entries = _RAND_4[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  entries_batch = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  dataout_width_cmp = _RAND_6[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  rls_entries = _RAND_7[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  h_bias_0_stride = _RAND_8[22:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  h_bias_1_stride = _RAND_9[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  slice_left = _RAND_10[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  is_winograd_d1 = _RAND_11[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  is_img_d1 = _RAND_12[33:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  data_bank = _RAND_13[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  datain_width = _RAND_14[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  datain_width_cmp = _RAND_15[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  datain_height_cmp = _RAND_16[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  datain_channel_cmp = _RAND_17[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  sub_h_total_g0 = _RAND_18[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  sub_h_total_g1 = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  sub_h_total_g2 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  sub_h_total_g3 = _RAND_21[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  sub_h_total_g4 = _RAND_22[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  sub_h_total_g5 = _RAND_23[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  sub_h_total_g6 = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  sub_h_total_g8 = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  sub_h_total_g9 = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  sub_h_total_g11 = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  sub_h_cmp_g0 = _RAND_28[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  sub_h_cmp_g1 = _RAND_29[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  conv_x_stride = _RAND_30[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  conv_y_stride = _RAND_31[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  batch_cmp = _RAND_32[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  pixel_x_init = _RAND_33[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  pixel_x_init_offset = _RAND_34[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  pixel_x_add = _RAND_35[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  pixel_x_byte_stride = _RAND_36[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  pixel_ch_stride = _RAND_37[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  x_dilate = _RAND_38[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  y_dilate = _RAND_39[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  pad_value = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  entries_cmp = _RAND_41[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  h_bias_2_stride = _RAND_42[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  h_bias_3_stride = _RAND_43[16:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  last_slices = _RAND_44[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  last_entries = _RAND_45[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  dat_entry_st = _RAND_46[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  dat_rsp_l3_pvld = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  dat_rsp_l1_pvld = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  dat_rsp_l0_pvld = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_1507 = _RAND_50[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_1501 = _RAND_51[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_1498 = _RAND_52[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_653 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_656 = _RAND_54[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_659 = _RAND_55[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_664 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_667 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_670 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_673 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_676 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_681 = _RAND_61[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_684 = _RAND_62[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_687 = _RAND_63[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_690 = _RAND_64[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_693 = _RAND_65[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_700 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_703 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_706 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_709 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_714 = _RAND_70[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_717 = _RAND_71[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_720 = _RAND_72[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_723 = _RAND_73[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  batch_cnt = _RAND_74[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  stripe_cnt = _RAND_75[6:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  sub_h_cnt = _RAND_76[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  dat_exec_valid_d1 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  dat_pipe_local_valid = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  dat_pipe_valid_d1 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  dat_req_bytes_d1 = _RAND_80[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  dataout_w_cnt = _RAND_81[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  dataout_w_ori = _RAND_82[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  datain_c_cnt = _RAND_83[10:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  datain_w_cnt = _RAND_84[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  datain_w_ori = _RAND_85[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  pixel_w_cnt = _RAND_86[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  pixel_w_ori = _RAND_87[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  pixel_w_ch_ori = _RAND_88[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  channel_op_cnt = _RAND_89[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  pixel_force_clr_d1 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  pixel_force_fetch_d1 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  datain_h_cnt = _RAND_92[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  datain_h_ori = _RAND_93[13:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  dat_req_valid_d1 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  dat_req_sub_w_d1 = _RAND_95[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  dat_req_sub_h_d1 = _RAND_96[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  dat_req_sub_c_d1 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  dat_req_ch_end_d1 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  dat_req_dummy_d1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  dat_req_cur_sub_h_d1 = _RAND_100[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  dat_req_sub_w_st_d1 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  dat_req_flag_d1 = _RAND_102[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  dat_req_rls_d1 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  c_bias = _RAND_104[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  c_bias_d1 = _RAND_105[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  h_bias_0_d1 = _RAND_106[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  h_bias_1_d1 = _RAND_107[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  h_bias_2_d1 = _RAND_108[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  h_bias_3_d1 = _RAND_109[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  w_bias_d1 = _RAND_110[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  dat_req_sub_h_addr_0 = _RAND_111[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  dat_req_sub_h_addr_1 = _RAND_112[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  dat_req_sub_h_addr_2 = _RAND_113[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  dat_req_sub_h_addr_3 = _RAND_114[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  sc2buf_dat_rd_en_out = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  sc2buf_dat_rd_addr_out = _RAND_116[18:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  dat_req_pipe_pvld = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  dat_req_exec_pvld = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  dat_req_exec_dummy = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  dat_req_pipe_sub_w = _RAND_120[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  dat_req_pipe_sub_h = _RAND_121[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  dat_req_pipe_sub_c = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  dat_req_pipe_ch_end = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  dat_req_pipe_bytes = _RAND_124[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  dat_req_pipe_dummy = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  dat_req_pipe_cur_sub_h = _RAND_126[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  dat_req_pipe_sub_w_st = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  dat_req_pipe_rls = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  dat_req_pipe_flag = _RAND_129[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_1276 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_1279 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_1282 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_1285 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_1288 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  dat_rsp_pipe_pvld = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_1295 = _RAND_136[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_1298 = _RAND_137[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_1301 = _RAND_138[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_1304 = _RAND_139[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_1307 = _RAND_140[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  dat_rsp_pipe_pd = _RAND_141[28:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_1314 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_1317 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_1320 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_1323 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_1326 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  dat_rsp_exec_pvld = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_1333 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_1336 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_1339 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_1342 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_1345 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  dat_rsp_exec_dummy = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_1352 = _RAND_154[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_1355 = _RAND_155[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_1358 = _RAND_156[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_1361 = _RAND_157[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_1364 = _RAND_158[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  dat_rsp_exec_sub_h = _RAND_159[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  dat_l0c0_dummy = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  dat_l1c0_dummy = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  dat_l2c0_dummy = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  dat_l3c0_dummy = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  dat_l0c1_dummy = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  dat_l1c1_dummy = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  dat_l2c1_dummy = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  dat_l3c1_dummy = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {16{`RANDOM}};
  dat_l0c0 = _RAND_168[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {16{`RANDOM}};
  dat_l1c0 = _RAND_169[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {16{`RANDOM}};
  dat_l2c0 = _RAND_170[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {16{`RANDOM}};
  dat_l3c0 = _RAND_171[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {16{`RANDOM}};
  dat_l0c1 = _RAND_172[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {16{`RANDOM}};
  dat_l1c1 = _RAND_173[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {16{`RANDOM}};
  dat_l2c1 = _RAND_174[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {16{`RANDOM}};
  dat_l3c1 = _RAND_175[511:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  rsp_sft_cnt_l0 = _RAND_176[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  rsp_sft_cnt_l1 = _RAND_177[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  rsp_sft_cnt_l2 = _RAND_178[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  rsp_sft_cnt_l3 = _RAND_179[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  rsp_sft_cnt_l0_ori = _RAND_180[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  rsp_sft_cnt_l1_ori = _RAND_181[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  rsp_sft_cnt_l2_ori = _RAND_182[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  rsp_sft_cnt_l3_ori = _RAND_183[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  dat_rsp_l2_pvld = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_1504 = _RAND_185[26:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {8{`RANDOM}};
  dat_rsp_l0_sft_d1 = _RAND_186[255:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {4{`RANDOM}};
  dat_rsp_l0_sft_d2 = _RAND_187[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {4{`RANDOM}};
  dat_rsp_l0_sft_d3 = _RAND_188[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {4{`RANDOM}};
  dat_rsp_l1_sft_d2 = _RAND_189[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {4{`RANDOM}};
  dat_rsp_l1_sft_d3 = _RAND_190[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {4{`RANDOM}};
  dat_rsp_l2_sft_d3 = _RAND_191[127:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  dat_out_pvld = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  dat_out_flag = _RAND_193[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  dat_out_bypass_mask_0 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  dat_out_bypass_mask_1 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  dat_out_bypass_mask_2 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  dat_out_bypass_mask_3 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  dat_out_bypass_mask_4 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  dat_out_bypass_mask_5 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  dat_out_bypass_mask_6 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  dat_out_bypass_mask_7 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  dat_out_bypass_mask_8 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  dat_out_bypass_mask_9 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  dat_out_bypass_mask_10 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  dat_out_bypass_mask_11 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  dat_out_bypass_mask_12 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  dat_out_bypass_mask_13 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  dat_out_bypass_mask_14 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  dat_out_bypass_mask_15 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  dat_out_bypass_mask_16 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  dat_out_bypass_mask_17 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  dat_out_bypass_mask_18 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  dat_out_bypass_mask_19 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  dat_out_bypass_mask_20 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  dat_out_bypass_mask_21 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  dat_out_bypass_mask_22 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  dat_out_bypass_mask_23 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  dat_out_bypass_mask_24 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  dat_out_bypass_mask_25 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  dat_out_bypass_mask_26 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  dat_out_bypass_mask_27 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  dat_out_bypass_mask_28 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  dat_out_bypass_mask_29 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  dat_out_bypass_mask_30 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  dat_out_bypass_mask_31 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  dat_out_bypass_mask_32 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  dat_out_bypass_mask_33 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  dat_out_bypass_mask_34 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  dat_out_bypass_mask_35 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  dat_out_bypass_mask_36 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  dat_out_bypass_mask_37 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  dat_out_bypass_mask_38 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  dat_out_bypass_mask_39 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  dat_out_bypass_mask_40 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  dat_out_bypass_mask_41 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  dat_out_bypass_mask_42 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  dat_out_bypass_mask_43 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  dat_out_bypass_mask_44 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  dat_out_bypass_mask_45 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  dat_out_bypass_mask_46 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  dat_out_bypass_mask_47 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  dat_out_bypass_mask_48 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  dat_out_bypass_mask_49 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  dat_out_bypass_mask_50 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  dat_out_bypass_mask_51 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  dat_out_bypass_mask_52 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  dat_out_bypass_mask_53 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  dat_out_bypass_mask_54 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  dat_out_bypass_mask_55 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  dat_out_bypass_mask_56 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  dat_out_bypass_mask_57 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  dat_out_bypass_mask_58 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  dat_out_bypass_mask_59 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  dat_out_bypass_mask_60 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  dat_out_bypass_mask_61 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  dat_out_bypass_mask_62 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  dat_out_bypass_mask_63 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  dat_out_bypass_data_0 = _RAND_258[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  dat_out_bypass_data_1 = _RAND_259[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  dat_out_bypass_data_2 = _RAND_260[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  dat_out_bypass_data_3 = _RAND_261[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  dat_out_bypass_data_4 = _RAND_262[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  dat_out_bypass_data_5 = _RAND_263[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  dat_out_bypass_data_6 = _RAND_264[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  dat_out_bypass_data_7 = _RAND_265[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  dat_out_bypass_data_8 = _RAND_266[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  dat_out_bypass_data_9 = _RAND_267[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  dat_out_bypass_data_10 = _RAND_268[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  dat_out_bypass_data_11 = _RAND_269[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  dat_out_bypass_data_12 = _RAND_270[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  dat_out_bypass_data_13 = _RAND_271[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  dat_out_bypass_data_14 = _RAND_272[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  dat_out_bypass_data_15 = _RAND_273[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  dat_out_bypass_data_16 = _RAND_274[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  dat_out_bypass_data_17 = _RAND_275[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  dat_out_bypass_data_18 = _RAND_276[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  dat_out_bypass_data_19 = _RAND_277[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  dat_out_bypass_data_20 = _RAND_278[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  dat_out_bypass_data_21 = _RAND_279[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  dat_out_bypass_data_22 = _RAND_280[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  dat_out_bypass_data_23 = _RAND_281[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  dat_out_bypass_data_24 = _RAND_282[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  dat_out_bypass_data_25 = _RAND_283[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  dat_out_bypass_data_26 = _RAND_284[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  dat_out_bypass_data_27 = _RAND_285[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  dat_out_bypass_data_28 = _RAND_286[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  dat_out_bypass_data_29 = _RAND_287[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  dat_out_bypass_data_30 = _RAND_288[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  dat_out_bypass_data_31 = _RAND_289[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  dat_out_bypass_data_32 = _RAND_290[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  dat_out_bypass_data_33 = _RAND_291[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  dat_out_bypass_data_34 = _RAND_292[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  dat_out_bypass_data_35 = _RAND_293[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  dat_out_bypass_data_36 = _RAND_294[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  dat_out_bypass_data_37 = _RAND_295[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  dat_out_bypass_data_38 = _RAND_296[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  dat_out_bypass_data_39 = _RAND_297[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  dat_out_bypass_data_40 = _RAND_298[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  dat_out_bypass_data_41 = _RAND_299[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  dat_out_bypass_data_42 = _RAND_300[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  dat_out_bypass_data_43 = _RAND_301[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  dat_out_bypass_data_44 = _RAND_302[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  dat_out_bypass_data_45 = _RAND_303[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  dat_out_bypass_data_46 = _RAND_304[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  dat_out_bypass_data_47 = _RAND_305[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  dat_out_bypass_data_48 = _RAND_306[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  dat_out_bypass_data_49 = _RAND_307[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  dat_out_bypass_data_50 = _RAND_308[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  dat_out_bypass_data_51 = _RAND_309[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  dat_out_bypass_data_52 = _RAND_310[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  dat_out_bypass_data_53 = _RAND_311[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  dat_out_bypass_data_54 = _RAND_312[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  dat_out_bypass_data_55 = _RAND_313[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  dat_out_bypass_data_56 = _RAND_314[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  dat_out_bypass_data_57 = _RAND_315[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  dat_out_bypass_data_58 = _RAND_316[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  dat_out_bypass_data_59 = _RAND_317[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  dat_out_bypass_data_60 = _RAND_318[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  dat_out_bypass_data_61 = _RAND_319[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  dat_out_bypass_data_62 = _RAND_320[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  dat_out_bypass_data_63 = _RAND_321[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_3147 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_3150 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_3153 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_3156 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_3159 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_3164 = _RAND_327[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_3167 = _RAND_328[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_3170 = _RAND_329[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_3173 = _RAND_330[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_3176 = _RAND_331[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  dl_out_pvld = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  dl_out_mask_0 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  dl_out_mask_1 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  dl_out_mask_2 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  dl_out_mask_3 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  dl_out_mask_4 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  dl_out_mask_5 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  dl_out_mask_6 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  dl_out_mask_7 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  dl_out_mask_8 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  dl_out_mask_9 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  dl_out_mask_10 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  dl_out_mask_11 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  dl_out_mask_12 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  dl_out_mask_13 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  dl_out_mask_14 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  dl_out_mask_15 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  dl_out_mask_16 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  dl_out_mask_17 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  dl_out_mask_18 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  dl_out_mask_19 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  dl_out_mask_20 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  dl_out_mask_21 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  dl_out_mask_22 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  dl_out_mask_23 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  dl_out_mask_24 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  dl_out_mask_25 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  dl_out_mask_26 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  dl_out_mask_27 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  dl_out_mask_28 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  dl_out_mask_29 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  dl_out_mask_30 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  dl_out_mask_31 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  dl_out_mask_32 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  dl_out_mask_33 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  dl_out_mask_34 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  dl_out_mask_35 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  dl_out_mask_36 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  dl_out_mask_37 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  dl_out_mask_38 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  dl_out_mask_39 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  dl_out_mask_40 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  dl_out_mask_41 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  dl_out_mask_42 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  dl_out_mask_43 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  dl_out_mask_44 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  dl_out_mask_45 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  dl_out_mask_46 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  dl_out_mask_47 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  dl_out_mask_48 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  dl_out_mask_49 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  dl_out_mask_50 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  dl_out_mask_51 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  dl_out_mask_52 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  dl_out_mask_53 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  dl_out_mask_54 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  dl_out_mask_55 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  dl_out_mask_56 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  dl_out_mask_57 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  dl_out_mask_58 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  dl_out_mask_59 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  dl_out_mask_60 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  dl_out_mask_61 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  dl_out_mask_62 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  dl_out_mask_63 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  dl_out_flag = _RAND_397[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  dl_out_data_0 = _RAND_398[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  dl_out_data_1 = _RAND_399[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  dl_out_data_2 = _RAND_400[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  dl_out_data_3 = _RAND_401[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  dl_out_data_4 = _RAND_402[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  dl_out_data_5 = _RAND_403[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  dl_out_data_6 = _RAND_404[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  dl_out_data_7 = _RAND_405[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  dl_out_data_8 = _RAND_406[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  dl_out_data_9 = _RAND_407[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  dl_out_data_10 = _RAND_408[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  dl_out_data_11 = _RAND_409[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  dl_out_data_12 = _RAND_410[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  dl_out_data_13 = _RAND_411[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  dl_out_data_14 = _RAND_412[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  dl_out_data_15 = _RAND_413[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  dl_out_data_16 = _RAND_414[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  dl_out_data_17 = _RAND_415[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  dl_out_data_18 = _RAND_416[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  dl_out_data_19 = _RAND_417[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  dl_out_data_20 = _RAND_418[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  dl_out_data_21 = _RAND_419[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  dl_out_data_22 = _RAND_420[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  dl_out_data_23 = _RAND_421[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  dl_out_data_24 = _RAND_422[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  dl_out_data_25 = _RAND_423[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  dl_out_data_26 = _RAND_424[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  dl_out_data_27 = _RAND_425[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  dl_out_data_28 = _RAND_426[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  dl_out_data_29 = _RAND_427[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  dl_out_data_30 = _RAND_428[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  dl_out_data_31 = _RAND_429[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  dl_out_data_32 = _RAND_430[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  dl_out_data_33 = _RAND_431[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  dl_out_data_34 = _RAND_432[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  dl_out_data_35 = _RAND_433[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  dl_out_data_36 = _RAND_434[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  dl_out_data_37 = _RAND_435[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  dl_out_data_38 = _RAND_436[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  dl_out_data_39 = _RAND_437[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  dl_out_data_40 = _RAND_438[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  dl_out_data_41 = _RAND_439[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  dl_out_data_42 = _RAND_440[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  dl_out_data_43 = _RAND_441[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  dl_out_data_44 = _RAND_442[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  dl_out_data_45 = _RAND_443[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  dl_out_data_46 = _RAND_444[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  dl_out_data_47 = _RAND_445[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  dl_out_data_48 = _RAND_446[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  dl_out_data_49 = _RAND_447[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  dl_out_data_50 = _RAND_448[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  dl_out_data_51 = _RAND_449[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  dl_out_data_52 = _RAND_450[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  dl_out_data_53 = _RAND_451[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  dl_out_data_54 = _RAND_452[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  dl_out_data_55 = _RAND_453[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  dl_out_data_56 = _RAND_454[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  dl_out_data_57 = _RAND_455[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  dl_out_data_58 = _RAND_456[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  dl_out_data_59 = _RAND_457[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  dl_out_data_60 = _RAND_458[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  dl_out_data_61 = _RAND_459[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  dl_out_data_62 = _RAND_460[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  dl_out_data_63 = _RAND_461[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  dl_out_pvld_d1 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_4582 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_4585 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_4589 = _RAND_465[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_4593 = _RAND_466[8:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_4861_0 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_4861_1 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_4861_2 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_4861_3 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_4861_4 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_4861_5 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_4861_6 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_4861_7 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_4861_8 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_4861_9 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_4861_10 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_4861_11 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_4861_12 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_4861_13 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_4861_14 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_4861_15 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_4861_16 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_4861_17 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_4861_18 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_4861_19 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_4861_20 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_4861_21 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_4861_22 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_4861_23 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_4861_24 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_4861_25 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_4861_26 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_4861_27 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_4861_28 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_4861_29 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_4861_30 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_4861_31 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_4861_32 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_4861_33 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_4861_34 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_4861_35 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_4861_36 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_4861_37 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_4861_38 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_4861_39 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_4861_40 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_4861_41 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_4861_42 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_4861_43 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_4861_44 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_4861_45 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_4861_46 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_4861_47 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_4861_48 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_4861_49 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_4861_50 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_4861_51 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_4861_52 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_4861_53 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_4861_54 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_4861_55 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_4861_56 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_4861_57 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_4861_58 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_4861_59 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_4861_60 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_4861_61 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_4861_62 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_4861_63 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_5388_0 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_5388_1 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_5388_2 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_5388_3 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_5388_4 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_5388_5 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_5388_6 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_5388_7 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_5388_8 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_5388_9 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_5388_10 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_5388_11 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_5388_12 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_5388_13 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_5388_14 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_5388_15 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_5388_16 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_5388_17 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_5388_18 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_5388_19 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_5388_20 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_5388_21 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_5388_22 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_5388_23 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_5388_24 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_5388_25 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_5388_26 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_5388_27 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_5388_28 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_5388_29 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_5388_30 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_5388_31 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_5388_32 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_5388_33 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_5388_34 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_5388_35 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_5388_36 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_5388_37 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_5388_38 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_5388_39 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_5388_40 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_5388_41 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_5388_42 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_5388_43 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_5388_44 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_5388_45 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_5388_46 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_5388_47 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_5388_48 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_5388_49 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_5388_50 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_5388_51 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_5388_52 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_5388_53 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_5388_54 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_5388_55 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_5388_56 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_5388_57 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_5388_58 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_5388_59 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_5388_60 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_5388_61 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_5388_62 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_5388_63 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_5649 = _RAND_595[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_5651 = _RAND_596[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_5653 = _RAND_597[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_5655 = _RAND_598[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_5657 = _RAND_599[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_5659 = _RAND_600[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_5661 = _RAND_601[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_5663 = _RAND_602[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_5665 = _RAND_603[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_5667 = _RAND_604[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_5669 = _RAND_605[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_5671 = _RAND_606[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_5673 = _RAND_607[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_5675 = _RAND_608[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_5677 = _RAND_609[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_5679 = _RAND_610[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_5681 = _RAND_611[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_5683 = _RAND_612[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_5685 = _RAND_613[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_5687 = _RAND_614[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_5689 = _RAND_615[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_5691 = _RAND_616[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_5693 = _RAND_617[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_5695 = _RAND_618[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_5697 = _RAND_619[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_5699 = _RAND_620[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_5701 = _RAND_621[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_5703 = _RAND_622[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_5705 = _RAND_623[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_5707 = _RAND_624[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_5709 = _RAND_625[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_5711 = _RAND_626[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_5713 = _RAND_627[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_5715 = _RAND_628[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_5717 = _RAND_629[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_5719 = _RAND_630[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_5721 = _RAND_631[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_5723 = _RAND_632[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_5725 = _RAND_633[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_5727 = _RAND_634[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_5729 = _RAND_635[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_5731 = _RAND_636[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_5733 = _RAND_637[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_5735 = _RAND_638[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_5737 = _RAND_639[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_5739 = _RAND_640[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_5741 = _RAND_641[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_5743 = _RAND_642[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_5745 = _RAND_643[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_5747 = _RAND_644[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_5749 = _RAND_645[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_5751 = _RAND_646[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_5753 = _RAND_647[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_5755 = _RAND_648[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_5757 = _RAND_649[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_5759 = _RAND_650[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_5761 = _RAND_651[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_5763 = _RAND_652[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_5765 = _RAND_653[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_5767 = _RAND_654[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_5769 = _RAND_655[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_5771 = _RAND_656[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_5773 = _RAND_657[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_5775 = _RAND_658[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_5777 = _RAND_659[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_5779 = _RAND_660[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_5781 = _RAND_661[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_5783 = _RAND_662[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_5785 = _RAND_663[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_5787 = _RAND_664[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_5789 = _RAND_665[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_5791 = _RAND_666[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_5793 = _RAND_667[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_5795 = _RAND_668[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_5797 = _RAND_669[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_5799 = _RAND_670[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_5801 = _RAND_671[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_5803 = _RAND_672[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_5805 = _RAND_673[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_5807 = _RAND_674[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_5809 = _RAND_675[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_5811 = _RAND_676[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_5813 = _RAND_677[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_5815 = _RAND_678[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_5817 = _RAND_679[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_5819 = _RAND_680[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_5821 = _RAND_681[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_5823 = _RAND_682[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_5825 = _RAND_683[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_5827 = _RAND_684[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_5829 = _RAND_685[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_5831 = _RAND_686[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_5833 = _RAND_687[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_5835 = _RAND_688[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_5837 = _RAND_689[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_5839 = _RAND_690[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_5841 = _RAND_691[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_5843 = _RAND_692[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_5845 = _RAND_693[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_5847 = _RAND_694[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_5849 = _RAND_695[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_5851 = _RAND_696[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_5853 = _RAND_697[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_5855 = _RAND_698[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_5857 = _RAND_699[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_5859 = _RAND_700[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_5861 = _RAND_701[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_5863 = _RAND_702[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_5865 = _RAND_703[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_5867 = _RAND_704[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_5869 = _RAND_705[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_5871 = _RAND_706[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_5873 = _RAND_707[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_5875 = _RAND_708[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_5877 = _RAND_709[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_5879 = _RAND_710[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_5881 = _RAND_711[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_5883 = _RAND_712[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_5885 = _RAND_713[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_5887 = _RAND_714[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_5889 = _RAND_715[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_5891 = _RAND_716[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_5893 = _RAND_717[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_5895 = _RAND_718[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_5897 = _RAND_719[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_5899 = _RAND_720[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_5901 = _RAND_721[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_5903 = _RAND_722[7:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge io_nvdla_core_clk) begin
    if (_T_207) begin
      layer_st_d1 <= 1'h0;
    end else begin
      layer_st_d1 <= layer_st;
    end
    if (_T_207) begin
      data_batch <= 6'h0;
    end else begin
      if (layer_st) begin
        data_batch <= 6'h1;
      end
    end
    if (_T_207) begin
      rls_slices <= 14'h0;
    end else begin
      if (layer_st) begin
        rls_slices <= {{1'd0}, rls_slices_w};
      end
    end
    if (_T_207) begin
      h_offset_slice <= 14'h0;
    end else begin
      if (layer_st) begin
        h_offset_slice <= {{2'd0}, h_offset_slice_w};
      end
    end
    if (_T_207) begin
      entries <= 17'h0;
    end else begin
      if (layer_st) begin
        entries <= entries_w;
      end
    end
    if (_T_207) begin
      entries_batch <= 15'h0;
    end else begin
      if (layer_st) begin
        entries_batch <= entries_batch_w;
      end
    end
    if (_T_207) begin
      dataout_width_cmp <= 13'h0;
    end else begin
      if (layer_st) begin
        dataout_width_cmp <= io_reg2dp_dataout_width;
      end
    end
    if (_T_207) begin
      rls_entries <= 29'h0;
    end else begin
      if (layer_st_d1) begin
        rls_entries <= slice_entries_w;
      end
    end
    if (_T_207) begin
      h_bias_0_stride <= 23'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_0_stride <= h_bias_0_stride_w;
      end
    end
    if (_T_207) begin
      h_bias_1_stride <= 31'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_1_stride <= h_bias_1_stride_w;
      end
    end
    if (_T_207) begin
      slice_left <= 14'h0;
    end else begin
      if (layer_st) begin
        if (io_reg2dp_skip_data_rls) begin
          slice_left <= _T_360;
        end else begin
          slice_left <= _T_362;
        end
      end
    end
    if (_T_207) begin
      is_winograd_d1 <= 22'h0;
    end else begin
      if (layer_st) begin
        is_winograd_d1 <= 22'h0;
      end
    end
    if (_T_207) begin
      is_img_d1 <= 34'h0;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          is_img_d1 <= 34'h3ffffffff;
        end else begin
          is_img_d1 <= 34'h0;
        end
      end
    end
    if (_T_207) begin
      data_bank <= 6'h0;
    end else begin
      if (layer_st) begin
        data_bank <= _T_549;
      end
    end
    if (_T_207) begin
      datain_width <= 14'h0;
    end else begin
      if (layer_st) begin
        datain_width <= _T_554;
      end
    end
    if (_T_207) begin
      datain_width_cmp <= 13'h0;
    end else begin
      if (layer_st) begin
        datain_width_cmp <= io_reg2dp_datain_width_ext;
      end
    end
    if (_T_207) begin
      datain_height_cmp <= 13'h0;
    end else begin
      if (layer_st) begin
        datain_height_cmp <= io_reg2dp_datain_height_ext;
      end
    end
    if (_T_207) begin
      datain_channel_cmp <= 11'h0;
    end else begin
      if (layer_st) begin
        datain_channel_cmp <= _T_558;
      end
    end
    if (_T_207) begin
      sub_h_total_g0 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g0 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g1 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g1 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g2 <= 2'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g2 <= _T_559;
      end
    end
    if (_T_207) begin
      sub_h_total_g3 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g3 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g4 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g4 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g5 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g5 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g6 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g6 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g8 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g8 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g9 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g9 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_total_g11 <= 3'h1;
    end else begin
      if (layer_st) begin
        sub_h_total_g11 <= sub_h_total_w;
      end
    end
    if (_T_207) begin
      sub_h_cmp_g0 <= 3'h1;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          sub_h_cmp_g0 <= sub_h_total_w;
        end else begin
          sub_h_cmp_g0 <= 3'h1;
        end
      end
    end
    if (_T_207) begin
      sub_h_cmp_g1 <= 3'h1;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          sub_h_cmp_g1 <= sub_h_total_w;
        end else begin
          sub_h_cmp_g1 <= 3'h1;
        end
      end
    end
    if (_T_207) begin
      conv_x_stride <= 4'h0;
    end else begin
      if (layer_st) begin
        conv_x_stride <= conv_x_stride_w;
      end
    end
    if (_T_207) begin
      conv_y_stride <= 4'h0;
    end else begin
      if (layer_st) begin
        conv_y_stride <= conv_y_stride_w;
      end
    end
    if (_T_207) begin
      batch_cmp <= 5'h0;
    end else begin
      if (layer_st) begin
        batch_cmp <= 5'h0;
      end
    end
    if (_T_207) begin
      pixel_x_init <= 7'h0;
    end else begin
      if (layer_st) begin
        if (_T_259) begin
          pixel_x_init <= _T_252;
        end else begin
          pixel_x_init <= {{1'd0}, _T_258};
        end
      end
    end
    if (_T_207) begin
      pixel_x_init_offset <= 7'h0;
    end else begin
      if (layer_st) begin
        pixel_x_init_offset <= pixel_x_init_offset_w;
      end
    end
    if (_T_207) begin
      pixel_x_add <= 8'h0;
    end else begin
      if (layer_st) begin
        if (_T_259) begin
          pixel_x_add <= _T_264;
        end else begin
          pixel_x_add <= {{1'd0}, _T_269};
        end
      end
    end
    if (_T_207) begin
      pixel_x_byte_stride <= 7'h0;
    end else begin
      if (layer_st) begin
        pixel_x_byte_stride <= {{1'd0}, pixel_x_stride_w};
      end
    end
    if (_T_207) begin
      pixel_ch_stride <= 12'h0;
    end else begin
      if (layer_st) begin
        pixel_ch_stride <= pixel_ch_stride_w;
      end
    end
    if (_T_207) begin
      x_dilate <= 6'h0;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          x_dilate <= 6'h1;
        end else begin
          x_dilate <= _T_278;
        end
      end
    end
    if (_T_207) begin
      y_dilate <= 6'h0;
    end else begin
      if (layer_st) begin
        if (is_img) begin
          y_dilate <= 6'h1;
        end else begin
          y_dilate <= _T_282;
        end
      end
    end
    if (_T_207) begin
      pad_value <= 16'h0;
    end else begin
      if (layer_st) begin
        pad_value <= io_reg2dp_pad_value;
      end
    end
    if (_T_207) begin
      entries_cmp <= 15'h0;
    end else begin
      if (layer_st) begin
        entries_cmp <= _T_562;
      end
    end
    if (_T_207) begin
      h_bias_2_stride <= 17'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_2_stride <= entries;
      end
    end
    if (_T_207) begin
      h_bias_3_stride <= 17'h0;
    end else begin
      if (layer_st_d1) begin
        h_bias_3_stride <= entries;
      end
    end
    if (_T_207) begin
      last_slices <= 14'h0;
    end else begin
      if (is_sg_done) begin
        last_slices <= slice_left;
      end
    end
    if (_T_207) begin
      last_entries <= 29'h0;
    end else begin
      if (is_sg_done) begin
        last_entries <= slice_entries_w;
      end
    end
    if (_T_207) begin
      dat_rsp_l3_pvld <= 1'h0;
    end else begin
      dat_rsp_l3_pvld <= dat_rsp_l2_pvld;
    end
    if (_T_207) begin
      dat_rsp_l1_pvld <= 1'h0;
    end else begin
      dat_rsp_l1_pvld <= dat_rsp_l0_pvld;
    end
    if (_T_207) begin
      dat_rsp_l0_pvld <= 1'h0;
    end else begin
      dat_rsp_l0_pvld <= dat_rsp_pipe_pvld;
    end
    if (_T_207) begin
      _T_1507 <= 27'h0;
    end else begin
      if (dat_rsp_l2_pvld) begin
        _T_1507 <= _T_1504;
      end
    end
    if (_T_207) begin
      _T_1501 <= 27'h0;
    end else begin
      if (dat_rsp_l0_pvld) begin
        _T_1501 <= _T_1498;
      end
    end
    if (_T_207) begin
      _T_1498 <= 27'h0;
    end else begin
      if (dat_rsp_pipe_pvld) begin
        _T_1498 <= _T_1516;
      end
    end
    if (_T_207) begin
      _T_653 <= 1'h0;
    end else begin
      _T_653 <= dat_rls;
    end
    if (_T_207) begin
      _T_656 <= 14'h0;
    end else begin
      if (dat_rls) begin
        if (sub_rls) begin
          _T_656 <= rls_slices;
        end else begin
          _T_656 <= last_slices;
        end
      end
    end
    if (_T_207) begin
      _T_659 <= 15'h0;
    end else begin
      if (dat_rls) begin
        _T_659 <= sc2cdma_dat_entries_w;
      end
    end
    if (_T_207) begin
      _T_664 <= 1'h0;
    end else begin
      _T_664 <= io_sg2dl_pd_valid;
    end
    if (_T_207) begin
      _T_667 <= 1'h0;
    end else begin
      _T_667 <= _T_664;
    end
    if (_T_207) begin
      _T_670 <= 1'h0;
    end else begin
      _T_670 <= _T_667;
    end
    if (_T_207) begin
      _T_673 <= 1'h0;
    end else begin
      _T_673 <= _T_670;
    end
    if (_T_207) begin
      _T_676 <= 1'h0;
    end else begin
      _T_676 <= _T_673;
    end
    if (_T_207) begin
      _T_681 <= 31'h0;
    end else begin
      if (io_sg2dl_pd_valid) begin
        _T_681 <= io_sg2dl_pd_bits;
      end
    end
    if (_T_207) begin
      _T_684 <= 31'h0;
    end else begin
      if (_T_664) begin
        _T_684 <= _T_681;
      end
    end
    if (_T_207) begin
      _T_687 <= 31'h0;
    end else begin
      if (_T_667) begin
        _T_687 <= _T_684;
      end
    end
    if (_T_207) begin
      _T_690 <= 31'h0;
    end else begin
      if (_T_670) begin
        _T_690 <= _T_687;
      end
    end
    if (_T_207) begin
      _T_693 <= 31'h0;
    end else begin
      if (_T_673) begin
        _T_693 <= _T_690;
      end
    end
    if (_T_207) begin
      _T_700 <= 1'h0;
    end else begin
      if (_T_694) begin
        _T_700 <= io_sg2dl_pd_valid;
      end else begin
        _T_700 <= _T_676;
      end
    end
    if (_T_207) begin
      _T_703 <= 1'h0;
    end else begin
      _T_703 <= _T_700;
    end
    if (_T_207) begin
      _T_706 <= 1'h0;
    end else begin
      _T_706 <= _T_703;
    end
    if (_T_207) begin
      _T_709 <= 1'h0;
    end else begin
      _T_709 <= _T_706;
    end
    if (_T_207) begin
      _T_714 <= 31'h0;
    end else begin
      if (dl_in_pvld) begin
        if (_T_695) begin
          _T_714 <= io_sg2dl_pd_bits;
        end else begin
          _T_714 <= _T_693;
        end
      end
    end
    if (_T_207) begin
      _T_717 <= 31'h0;
    end else begin
      if (_T_700) begin
        _T_717 <= _T_714;
      end
    end
    if (_T_207) begin
      _T_720 <= 31'h0;
    end else begin
      if (_T_703) begin
        _T_720 <= _T_717;
      end
    end
    if (_T_207) begin
      _T_723 <= 31'h0;
    end else begin
      if (_T_706) begin
        _T_723 <= _T_720;
      end
    end
    if (_T_207) begin
      batch_cnt <= 5'h0;
    end else begin
      batch_cnt <= _GEN_68[4:0];
    end
    if (_T_207) begin
      stripe_cnt <= 7'h0;
    end else begin
      if (stripe_cnt_reg_en) begin
        if (layer_st) begin
          stripe_cnt <= 7'h0;
        end else begin
          if (!(_T_787)) begin
            if (is_stripe_end) begin
              stripe_cnt <= 7'h0;
            end else begin
              stripe_cnt <= stripe_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_207) begin
      sub_h_cnt <= 2'h0;
    end else begin
      sub_h_cnt <= _GEN_69[1:0];
    end
    if (_T_207) begin
      dat_exec_valid_d1 <= 1'h0;
    end else begin
      if (dl_pvld) begin
        dat_exec_valid_d1 <= 1'h1;
      end else begin
        if (_T_815) begin
          dat_exec_valid_d1 <= 1'h0;
        end
      end
    end
    if (_T_207) begin
      dat_pipe_local_valid <= 1'h0;
    end else begin
      if (_T_799) begin
        dat_pipe_local_valid <= 1'h0;
      end else begin
        if (dl_pvld) begin
          dat_pipe_local_valid <= 1'h1;
        end
      end
    end
    if (_T_207) begin
      dat_pipe_valid_d1 <= 1'h0;
    end else begin
      dat_pipe_valid_d1 <= dat_pipe_valid;
    end
    if (_T_207) begin
      dat_req_bytes_d1 <= 8'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_bytes_d1 <= dat_req_bytes;
      end
    end
    if (_T_207) begin
      dataout_w_cnt <= 13'h0;
    end else begin
      if (dataout_w_cnt_reg_en) begin
        if (layer_st) begin
          dataout_w_cnt <= {{9'd0}, dataout_w_init};
        end else begin
          if (_T_831) begin
            dataout_w_cnt <= dataout_w_ori;
          end else begin
            if (is_w_end) begin
              dataout_w_cnt <= {{9'd0}, dataout_w_init};
            end else begin
              dataout_w_cnt <= dataout_w_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_207) begin
      dataout_w_ori <= 13'h0;
    end else begin
      if (dataout_w_ori_reg_en) begin
        if (layer_st) begin
          dataout_w_ori <= {{9'd0}, dataout_w_init};
        end else begin
          if (!(_T_831)) begin
            if (is_w_end) begin
              dataout_w_ori <= {{9'd0}, dataout_w_init};
            end else begin
              dataout_w_ori <= dataout_w_cnt_inc;
            end
          end
        end
      end
    end
    if (_T_207) begin
      datain_c_cnt <= 11'h0;
    end else begin
      if (datain_c_cnt_reg_en) begin
        if (layer_st) begin
          datain_c_cnt <= 11'h0;
        end else begin
          if (dl_channel_end) begin
            datain_c_cnt <= 11'h0;
          end else begin
            datain_c_cnt <= _T_846;
          end
        end
      end
    end
    if (_T_207) begin
      datain_w_cnt <= 14'h0;
    end else begin
      datain_w_cnt <= _GEN_75[13:0];
    end
    if (_T_207) begin
      datain_w_ori <= 14'h0;
    end else begin
      datain_w_ori <= _GEN_77[13:0];
    end
    if (_T_207) begin
      pixel_w_cnt <= 16'h0;
    end else begin
      pixel_w_cnt <= _GEN_76[15:0];
    end
    if (_T_207) begin
      pixel_w_ori <= 16'h0;
    end else begin
      pixel_w_ori <= _GEN_78[15:0];
    end
    if (_T_207) begin
      pixel_w_ch_ori <= 16'h0;
    end else begin
      pixel_w_ch_ori <= _GEN_79[15:0];
    end
    if (_T_207) begin
      channel_op_cnt <= 13'h2;
    end else begin
      channel_op_cnt <= _T_905[12:0];
    end
    if (_T_207) begin
      pixel_force_clr_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        pixel_force_clr_d1 <= pixel_force_clr;
      end
    end
    if (_T_207) begin
      pixel_force_fetch_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        if (_T_950) begin
          pixel_force_fetch_d1 <= 1'h1;
        end else begin
          if (pixel_force_clr_d1) begin
            pixel_force_fetch_d1 <= 1'h0;
          end
        end
      end
    end
    if (_T_207) begin
      datain_h_cnt <= 14'h0;
    end else begin
      datain_h_cnt <= _GEN_80[13:0];
    end
    if (_T_207) begin
      datain_h_ori <= 14'h0;
    end else begin
      datain_h_ori <= _GEN_81[13:0];
    end
    if (_T_207) begin
      dat_req_valid_d1 <= 1'h0;
    end else begin
      dat_req_valid_d1 <= dat_req_valid;
    end
    if (_T_207) begin
      dat_req_sub_w_d1 <= 2'h0;
    end else begin
      if (dat_exec_valid) begin
        if (_T_1011) begin
          dat_req_sub_w_d1 <= {{1'd0}, _T_1013};
        end else begin
          dat_req_sub_w_d1 <= _T_1014;
        end
      end
    end
    if (_T_207) begin
      dat_req_sub_h_d1 <= 2'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_sub_h_d1 <= sub_h_cnt;
      end
    end
    if (_T_207) begin
      dat_req_sub_c_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        if (_T_1009) begin
          dat_req_sub_c_d1 <= _T_1010;
        end else begin
          dat_req_sub_c_d1 <= dl_block_end;
        end
      end
    end
    if (_T_207) begin
      dat_req_ch_end_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_ch_end_d1 <= is_last_channel;
      end
    end
    if (_T_207) begin
      dat_req_dummy_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        if (_T_998) begin
          dat_req_dummy_d1 <= dat_img_req_dummy;
        end else begin
          if (_T_999) begin
            dat_req_dummy_d1 <= 1'h0;
          end else begin
            dat_req_dummy_d1 <= dat_conv_req_dummy;
          end
        end
      end
    end
    if (_T_207) begin
      dat_req_cur_sub_h_d1 <= 2'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_cur_sub_h_d1 <= dl_cur_sub_h;
      end
    end
    if (_T_207) begin
      dat_req_sub_w_st_d1 <= 1'h0;
    end else begin
      if (dat_req_sub_w_st_en) begin
        dat_req_sub_w_st_d1 <= dl_pvld;
      end
    end
    if (_T_207) begin
      dat_req_flag_d1 <= 9'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_flag_d1 <= dat_req_flag_w;
      end
    end
    if (_T_207) begin
      dat_req_rls_d1 <= 1'h0;
    end else begin
      if (dat_exec_valid) begin
        dat_req_rls_d1 <= _T_1041;
      end
    end
    if (_T_207) begin
      c_bias <= 13'h0;
    end else begin
      if (datain_c_cnt_reg_en) begin
        if (layer_st) begin
          c_bias <= 13'h0;
        end else begin
          if (_T_1061) begin
            c_bias <= 13'h0;
          end else begin
            c_bias <= _T_1064;
          end
        end
      end
    end
    if (_T_207) begin
      c_bias_d1 <= 13'h0;
    end else begin
      if (c_bias_d1_reg_en) begin
        c_bias_d1 <= c_bias;
      end
    end
    if (_T_207) begin
      h_bias_0_d1 <= 13'h0;
    end else begin
      if (_T_1101) begin
        h_bias_0_d1 <= h_bias_0_w;
      end
    end
    if (_T_207) begin
      h_bias_1_d1 <= 13'h0;
    end else begin
      if (_T_1101) begin
        h_bias_1_d1 <= h_bias_1_w;
      end
    end
    if (_T_207) begin
      h_bias_2_d1 <= 13'h0;
    end else begin
      if (_T_1101) begin
        h_bias_2_d1 <= h_bias_2_w;
      end
    end
    if (_T_207) begin
      h_bias_3_d1 <= 13'h0;
    end else begin
      if (_T_1102) begin
        h_bias_3_d1 <= h_bias_3_w;
      end
    end
    if (_T_207) begin
      w_bias_d1 <= 13'h0;
    end else begin
      w_bias_d1 <= _GEN_99[12:0];
    end
    if (_T_207) begin
      dat_req_sub_h_addr_0 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_0 <= _GEN_100[12:0];
    end
    if (_T_207) begin
      dat_req_sub_h_addr_1 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_1 <= _GEN_101[12:0];
    end
    if (_T_207) begin
      dat_req_sub_h_addr_2 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_2 <= _GEN_102[12:0];
    end
    if (_T_207) begin
      dat_req_sub_h_addr_3 <= 13'h1fff;
    end else begin
      dat_req_sub_h_addr_3 <= _GEN_103[12:0];
    end
    if (_T_207) begin
      sc2buf_dat_rd_en_out <= 1'h0;
    end else begin
      sc2buf_dat_rd_en_out <= sc2buf_dat_rd_en_w;
    end
    if (_T_207) begin
      sc2buf_dat_rd_addr_out <= 19'h1fff;
    end else begin
      if (_T_1261) begin
        if (_T_1215) begin
          sc2buf_dat_rd_addr_out <= 19'h1fff;
        end else begin
          if (is_dat_req_addr_wrap) begin
            sc2buf_dat_rd_addr_out <= dat_req_addr_wrap;
          end else begin
            sc2buf_dat_rd_addr_out <= {{1'd0}, dat_req_addr_sum};
          end
        end
      end
    end
    if (_T_207) begin
      dat_req_pipe_pvld <= 1'h0;
    end else begin
      dat_req_pipe_pvld <= dat_pipe_valid_d1;
    end
    if (_T_207) begin
      dat_req_exec_pvld <= 1'h0;
    end else begin
      dat_req_exec_pvld <= dat_exec_valid_d1;
    end
    if (_T_207) begin
      dat_req_exec_dummy <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_exec_dummy <= dat_req_dummy_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_sub_w <= 2'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_w <= dat_req_sub_w_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_sub_h <= 2'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_h <= dat_req_sub_h_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_sub_c <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_c <= dat_req_sub_c_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_ch_end <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_ch_end <= dat_req_ch_end_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_bytes <= 8'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_bytes <= dat_req_bytes_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_dummy <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_dummy <= dat_req_dummy_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_cur_sub_h <= 2'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_cur_sub_h <= dat_req_cur_sub_h_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_sub_w_st <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_sub_w_st <= dat_req_sub_w_st_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_rls <= 1'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_rls <= dat_req_rls_d1;
      end
    end
    if (_T_207) begin
      dat_req_pipe_flag <= 9'h0;
    end else begin
      if (dat_exec_valid_d1) begin
        dat_req_pipe_flag <= dat_req_flag_d1;
      end
    end
    if (_T_207) begin
      _T_1276 <= 1'h0;
    end else begin
      _T_1276 <= dat_req_pipe_pvld;
    end
    if (_T_207) begin
      _T_1279 <= 1'h0;
    end else begin
      _T_1279 <= _T_1276;
    end
    if (_T_207) begin
      _T_1282 <= 1'h0;
    end else begin
      _T_1282 <= _T_1279;
    end
    if (_T_207) begin
      _T_1285 <= 1'h0;
    end else begin
      _T_1285 <= _T_1282;
    end
    if (_T_207) begin
      _T_1288 <= 1'h0;
    end else begin
      _T_1288 <= _T_1285;
    end
    if (_T_207) begin
      dat_rsp_pipe_pvld <= 1'h0;
    end else begin
      dat_rsp_pipe_pvld <= _T_1288;
    end
    if (_T_207) begin
      _T_1295 <= 29'h0;
    end else begin
      if (dat_req_pipe_pvld) begin
        _T_1295 <= dat_req_pipe_pd;
      end
    end
    if (_T_207) begin
      _T_1298 <= 29'h0;
    end else begin
      if (_T_1276) begin
        _T_1298 <= _T_1295;
      end
    end
    if (_T_207) begin
      _T_1301 <= 29'h0;
    end else begin
      if (_T_1279) begin
        _T_1301 <= _T_1298;
      end
    end
    if (_T_207) begin
      _T_1304 <= 29'h0;
    end else begin
      if (_T_1282) begin
        _T_1304 <= _T_1301;
      end
    end
    if (_T_207) begin
      _T_1307 <= 29'h0;
    end else begin
      if (_T_1285) begin
        _T_1307 <= _T_1304;
      end
    end
    if (_T_207) begin
      dat_rsp_pipe_pd <= 29'h0;
    end else begin
      if (_T_1288) begin
        dat_rsp_pipe_pd <= _T_1307;
      end
    end
    if (_T_207) begin
      _T_1314 <= 1'h0;
    end else begin
      _T_1314 <= dat_req_exec_pvld;
    end
    if (_T_207) begin
      _T_1317 <= 1'h0;
    end else begin
      _T_1317 <= _T_1314;
    end
    if (_T_207) begin
      _T_1320 <= 1'h0;
    end else begin
      _T_1320 <= _T_1317;
    end
    if (_T_207) begin
      _T_1323 <= 1'h0;
    end else begin
      _T_1323 <= _T_1320;
    end
    if (_T_207) begin
      _T_1326 <= 1'h0;
    end else begin
      _T_1326 <= _T_1323;
    end
    if (_T_207) begin
      dat_rsp_exec_pvld <= 1'h0;
    end else begin
      dat_rsp_exec_pvld <= _T_1326;
    end
    if (_T_207) begin
      _T_1333 <= 1'h0;
    end else begin
      if (dat_req_exec_pvld) begin
        _T_1333 <= dat_req_exec_dummy;
      end
    end
    if (_T_207) begin
      _T_1336 <= 1'h0;
    end else begin
      if (_T_1314) begin
        _T_1336 <= _T_1333;
      end
    end
    if (_T_207) begin
      _T_1339 <= 1'h0;
    end else begin
      if (_T_1317) begin
        _T_1339 <= _T_1336;
      end
    end
    if (_T_207) begin
      _T_1342 <= 1'h0;
    end else begin
      if (_T_1320) begin
        _T_1342 <= _T_1339;
      end
    end
    if (_T_207) begin
      _T_1345 <= 1'h0;
    end else begin
      if (_T_1323) begin
        _T_1345 <= _T_1342;
      end
    end
    if (_T_207) begin
      dat_rsp_exec_dummy <= 1'h0;
    end else begin
      if (_T_1326) begin
        dat_rsp_exec_dummy <= _T_1345;
      end
    end
    if (_T_207) begin
      _T_1352 <= 2'h0;
    end else begin
      if (dat_req_exec_pvld) begin
        _T_1352 <= 2'h0;
      end
    end
    if (_T_207) begin
      _T_1355 <= 2'h0;
    end else begin
      if (_T_1314) begin
        _T_1355 <= _T_1352;
      end
    end
    if (_T_207) begin
      _T_1358 <= 2'h0;
    end else begin
      if (_T_1317) begin
        _T_1358 <= _T_1355;
      end
    end
    if (_T_207) begin
      _T_1361 <= 2'h0;
    end else begin
      if (_T_1320) begin
        _T_1361 <= _T_1358;
      end
    end
    if (_T_207) begin
      _T_1364 <= 2'h0;
    end else begin
      if (_T_1323) begin
        _T_1364 <= _T_1361;
      end
    end
    if (_T_207) begin
      dat_rsp_exec_sub_h <= 2'h0;
    end else begin
      if (_T_1326) begin
        dat_rsp_exec_sub_h <= _T_1364;
      end
    end
    if (_T_207) begin
      dat_l0c0_dummy <= 1'h1;
    end else begin
      if (dat_l0c0_en) begin
        dat_l0c0_dummy <= 1'h0;
      end else begin
        if (dat_dummy_l0_en) begin
          dat_l0c0_dummy <= 1'h1;
        end
      end
    end
    if (_T_207) begin
      dat_l1c0_dummy <= 1'h1;
    end else begin
      if (dat_l1c0_en) begin
        dat_l1c0_dummy <= 1'h0;
      end else begin
        if (dat_dummy_l1_en) begin
          dat_l1c0_dummy <= 1'h1;
        end
      end
    end
    if (_T_207) begin
      dat_l2c0_dummy <= 1'h1;
    end else begin
      if (dat_l2c0_en) begin
        dat_l2c0_dummy <= 1'h0;
      end else begin
        if (dat_dummy_l2_en) begin
          dat_l2c0_dummy <= 1'h1;
        end
      end
    end
    if (_T_207) begin
      dat_l3c0_dummy <= 1'h1;
    end else begin
      if (dat_l3c0_en) begin
        dat_l3c0_dummy <= 1'h0;
      end else begin
        if (dat_dummy_l3_en) begin
          dat_l3c0_dummy <= 1'h1;
        end
      end
    end
    if (_T_207) begin
      dat_l0c1_dummy <= 1'h1;
    end else begin
      if (dat_l0c1_en) begin
        dat_l0c1_dummy <= 1'h0;
      end else begin
        if (dat_l0_set) begin
          dat_l0c1_dummy <= dat_l0c0_dummy;
        end
      end
    end
    if (_T_207) begin
      dat_l1c1_dummy <= 1'h1;
    end else begin
      if (dat_l1c1_en) begin
        dat_l1c1_dummy <= 1'h0;
      end else begin
        if (_T_1455) begin
          dat_l1c1_dummy <= dat_l1c0_dummy;
        end
      end
    end
    if (_T_207) begin
      dat_l2c1_dummy <= 1'h1;
    end else begin
      if (dat_l2c1_en) begin
        dat_l2c1_dummy <= 1'h0;
      end else begin
        if (_T_1460) begin
          dat_l2c1_dummy <= dat_l2c0_dummy;
        end
      end
    end
    if (_T_207) begin
      dat_l3c1_dummy <= 1'h1;
    end else begin
      if (dat_l3c1_en) begin
        dat_l3c1_dummy <= 1'h0;
      end else begin
        if (_T_1465) begin
          dat_l3c1_dummy <= dat_l3c0_dummy;
        end
      end
    end
    if (dat_l0c0_en) begin
      dat_l0c0 <= io_sc2buf_dat_rd_data_bits;
    end
    if (dat_l1c0_en) begin
      dat_l1c0 <= io_sc2buf_dat_rd_data_bits;
    end
    if (dat_l2c0_en) begin
      dat_l2c0 <= io_sc2buf_dat_rd_data_bits;
    end
    if (dat_l3c0_en) begin
      dat_l3c0 <= io_sc2buf_dat_rd_data_bits;
    end
    if (dat_l0c1_en) begin
      dat_l0c1 <= dat_l0c0;
    end
    if (dat_l1c1_en) begin
      dat_l1c1 <= dat_l1c0;
    end
    if (dat_l2c1_en) begin
      dat_l2c1 <= dat_l2c0;
    end
    if (dat_l3c1_en) begin
      dat_l3c1 <= dat_l3c0;
    end
    if (_T_207) begin
      rsp_sft_cnt_l0 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l0_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l0 <= 8'h40;
        end else begin
          if (_T_1583) begin
            rsp_sft_cnt_l0 <= rsp_sft_cnt_l0_ori;
          end else begin
            if (_T_1584) begin
              rsp_sft_cnt_l0 <= 8'h40;
            end else begin
              if (dat_dummy_l0_en) begin
                rsp_sft_cnt_l0 <= _T_1587;
              end else begin
                rsp_sft_cnt_l0 <= rsp_sft_cnt_l0_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l1 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l1_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l1 <= 8'h40;
        end else begin
          if (_T_1593) begin
            rsp_sft_cnt_l1 <= rsp_sft_cnt_l1_ori;
          end else begin
            if (_T_1594) begin
              rsp_sft_cnt_l1 <= 8'h40;
            end else begin
              if (dat_dummy_l1_en) begin
                rsp_sft_cnt_l1 <= _T_1597;
              end else begin
                rsp_sft_cnt_l1 <= rsp_sft_cnt_l1_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l2 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l2_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l2 <= 8'h40;
        end else begin
          if (_T_1603) begin
            rsp_sft_cnt_l2 <= rsp_sft_cnt_l2_ori;
          end else begin
            if (_T_1604) begin
              rsp_sft_cnt_l2 <= 8'h40;
            end else begin
              if (dat_dummy_l2_en) begin
                rsp_sft_cnt_l2 <= _T_1607;
              end else begin
                rsp_sft_cnt_l2 <= rsp_sft_cnt_l2_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l3 <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l3_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l3 <= 8'h40;
        end else begin
          if (_T_1613) begin
            rsp_sft_cnt_l3 <= rsp_sft_cnt_l3_ori;
          end else begin
            if (_T_1614) begin
              rsp_sft_cnt_l3 <= 8'h40;
            end else begin
              if (dat_dummy_l3_en) begin
                rsp_sft_cnt_l3 <= _T_1617;
              end else begin
                rsp_sft_cnt_l3 <= rsp_sft_cnt_l3_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l0_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l0_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l0_ori <= 8'h40;
        end else begin
          if (!(_T_1583)) begin
            if (_T_1584) begin
              rsp_sft_cnt_l0_ori <= 8'h40;
            end else begin
              if (dat_dummy_l0_en) begin
                rsp_sft_cnt_l0_ori <= _T_1587;
              end else begin
                rsp_sft_cnt_l0_ori <= rsp_sft_cnt_l0_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l1_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l1_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l1_ori <= 8'h40;
        end else begin
          if (!(_T_1593)) begin
            if (_T_1594) begin
              rsp_sft_cnt_l1_ori <= 8'h40;
            end else begin
              if (dat_dummy_l1_en) begin
                rsp_sft_cnt_l1_ori <= _T_1597;
              end else begin
                rsp_sft_cnt_l1_ori <= rsp_sft_cnt_l1_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l2_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l2_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l2_ori <= 8'h40;
        end else begin
          if (!(_T_1603)) begin
            if (_T_1604) begin
              rsp_sft_cnt_l2_ori <= 8'h40;
            end else begin
              if (dat_dummy_l2_en) begin
                rsp_sft_cnt_l2_ori <= _T_1607;
              end else begin
                rsp_sft_cnt_l2_ori <= rsp_sft_cnt_l2_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      rsp_sft_cnt_l3_ori <= 8'h0;
    end else begin
      if (rsp_sft_cnt_l3_ori_en) begin
        if (layer_st) begin
          rsp_sft_cnt_l3_ori <= 8'h40;
        end else begin
          if (!(_T_1613)) begin
            if (_T_1614) begin
              rsp_sft_cnt_l3_ori <= 8'h40;
            end else begin
              if (dat_dummy_l3_en) begin
                rsp_sft_cnt_l3_ori <= _T_1617;
              end else begin
                rsp_sft_cnt_l3_ori <= rsp_sft_cnt_l3_inc;
              end
            end
          end
        end
      end
    end
    if (_T_207) begin
      dat_rsp_l2_pvld <= 1'h0;
    end else begin
      dat_rsp_l2_pvld <= dat_rsp_l1_pvld;
    end
    if (_T_207) begin
      _T_1504 <= 27'h0;
    end else begin
      if (dat_rsp_l1_pvld) begin
        _T_1504 <= _T_1501;
      end
    end
    dat_rsp_l0_sft_d1 <= _GEN_154[255:0];
    dat_rsp_l0_sft_d2 <= _GEN_155[127:0];
    if (dat_rsp_sft_d3_en) begin
      dat_rsp_l0_sft_d3 <= dat_rsp_l0_sft_d2;
    end
    dat_rsp_l1_sft_d2 <= _GEN_156[127:0];
    if (dat_rsp_sft_d3_en) begin
      dat_rsp_l1_sft_d3 <= dat_rsp_l1_sft_d2;
    end
    dat_rsp_l2_sft_d3 <= _GEN_159[127:0];
    if (_T_207) begin
      dat_out_pvld <= 1'h0;
    end else begin
      if (_T_3177) begin
        dat_out_pvld <= _T_3159;
      end else begin
        dat_out_pvld <= dat_rsp_pvld;
      end
    end
    if (_T_207) begin
      dat_out_flag <= 9'h0;
    end else begin
      if (dat_out_pvld_w) begin
        if (_T_3178) begin
          dat_out_flag <= _T_3176;
        end else begin
          dat_out_flag <= dat_rsp_flag;
        end
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_0 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_0 <= dat_rsp_mask_w_0;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_1 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_1 <= dat_rsp_mask_w_1;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_2 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_2 <= dat_rsp_mask_w_2;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_3 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_3 <= dat_rsp_mask_w_3;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_4 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_4 <= dat_rsp_mask_w_4;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_5 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_5 <= dat_rsp_mask_w_5;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_6 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_6 <= dat_rsp_mask_w_6;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_7 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_7 <= dat_rsp_mask_w_7;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_8 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_8 <= dat_rsp_mask_w_8;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_9 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_9 <= dat_rsp_mask_w_9;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_10 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_10 <= dat_rsp_mask_w_10;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_11 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_11 <= dat_rsp_mask_w_11;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_12 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_12 <= dat_rsp_mask_w_12;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_13 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_13 <= dat_rsp_mask_w_13;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_14 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_14 <= dat_rsp_mask_w_14;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_15 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_15 <= dat_rsp_mask_w_15;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_16 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_16 <= dat_rsp_mask_w_16;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_17 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_17 <= dat_rsp_mask_w_17;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_18 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_18 <= dat_rsp_mask_w_18;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_19 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_19 <= dat_rsp_mask_w_19;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_20 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_20 <= dat_rsp_mask_w_20;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_21 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_21 <= dat_rsp_mask_w_21;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_22 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_22 <= dat_rsp_mask_w_22;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_23 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_23 <= dat_rsp_mask_w_23;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_24 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_24 <= dat_rsp_mask_w_24;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_25 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_25 <= dat_rsp_mask_w_25;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_26 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_26 <= dat_rsp_mask_w_26;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_27 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_27 <= dat_rsp_mask_w_27;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_28 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_28 <= dat_rsp_mask_w_28;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_29 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_29 <= dat_rsp_mask_w_29;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_30 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_30 <= dat_rsp_mask_w_30;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_31 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_31 <= dat_rsp_mask_w_31;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_32 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_32 <= dat_rsp_mask_w_32;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_33 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_33 <= dat_rsp_mask_w_33;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_34 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_34 <= dat_rsp_mask_w_34;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_35 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_35 <= dat_rsp_mask_w_35;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_36 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_36 <= dat_rsp_mask_w_36;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_37 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_37 <= dat_rsp_mask_w_37;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_38 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_38 <= dat_rsp_mask_w_38;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_39 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_39 <= dat_rsp_mask_w_39;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_40 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_40 <= dat_rsp_mask_w_40;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_41 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_41 <= dat_rsp_mask_w_41;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_42 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_42 <= dat_rsp_mask_w_42;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_43 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_43 <= dat_rsp_mask_w_43;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_44 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_44 <= dat_rsp_mask_w_44;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_45 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_45 <= dat_rsp_mask_w_45;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_46 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_46 <= dat_rsp_mask_w_46;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_47 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_47 <= dat_rsp_mask_w_47;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_48 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_48 <= dat_rsp_mask_w_48;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_49 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_49 <= dat_rsp_mask_w_49;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_50 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_50 <= dat_rsp_mask_w_50;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_51 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_51 <= dat_rsp_mask_w_51;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_52 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_52 <= dat_rsp_mask_w_52;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_53 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_53 <= dat_rsp_mask_w_53;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_54 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_54 <= dat_rsp_mask_w_54;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_55 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_55 <= dat_rsp_mask_w_55;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_56 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_56 <= dat_rsp_mask_w_56;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_57 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_57 <= dat_rsp_mask_w_57;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_58 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_58 <= dat_rsp_mask_w_58;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_59 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_59 <= dat_rsp_mask_w_59;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_60 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_60 <= dat_rsp_mask_w_60;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_61 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_61 <= dat_rsp_mask_w_61;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_62 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_62 <= dat_rsp_mask_w_62;
      end
    end
    if (_T_207) begin
      dat_out_bypass_mask_63 <= 1'h0;
    end else begin
      if (dat_rsp_p0_vld_w) begin
        dat_out_bypass_mask_63 <= dat_rsp_mask_w_63;
      end
    end
    if (_T_3179) begin
      if (_T_2080) begin
        dat_out_bypass_data_0 <= dat_rsp_img_0;
      end else begin
        dat_out_bypass_data_0 <= dat_rsp_conv_0;
      end
    end
    if (_T_3180) begin
      if (_T_2080) begin
        dat_out_bypass_data_1 <= dat_rsp_img_1;
      end else begin
        dat_out_bypass_data_1 <= dat_rsp_conv_1;
      end
    end
    if (_T_3181) begin
      if (_T_2080) begin
        dat_out_bypass_data_2 <= dat_rsp_img_2;
      end else begin
        dat_out_bypass_data_2 <= dat_rsp_conv_2;
      end
    end
    if (_T_3182) begin
      if (_T_2080) begin
        dat_out_bypass_data_3 <= dat_rsp_img_3;
      end else begin
        dat_out_bypass_data_3 <= dat_rsp_conv_3;
      end
    end
    if (_T_3183) begin
      if (_T_2080) begin
        dat_out_bypass_data_4 <= dat_rsp_img_4;
      end else begin
        dat_out_bypass_data_4 <= dat_rsp_conv_4;
      end
    end
    if (_T_3184) begin
      if (_T_2080) begin
        dat_out_bypass_data_5 <= dat_rsp_img_5;
      end else begin
        dat_out_bypass_data_5 <= dat_rsp_conv_5;
      end
    end
    if (_T_3185) begin
      if (_T_2080) begin
        dat_out_bypass_data_6 <= dat_rsp_img_6;
      end else begin
        dat_out_bypass_data_6 <= dat_rsp_conv_6;
      end
    end
    if (_T_3186) begin
      if (_T_2080) begin
        dat_out_bypass_data_7 <= dat_rsp_img_7;
      end else begin
        dat_out_bypass_data_7 <= dat_rsp_conv_7;
      end
    end
    if (_T_3187) begin
      if (_T_2080) begin
        dat_out_bypass_data_8 <= dat_rsp_img_8;
      end else begin
        dat_out_bypass_data_8 <= dat_rsp_conv_8;
      end
    end
    if (_T_3188) begin
      if (_T_2080) begin
        dat_out_bypass_data_9 <= dat_rsp_img_9;
      end else begin
        dat_out_bypass_data_9 <= dat_rsp_conv_9;
      end
    end
    if (_T_3189) begin
      if (_T_2080) begin
        dat_out_bypass_data_10 <= dat_rsp_img_10;
      end else begin
        dat_out_bypass_data_10 <= dat_rsp_conv_10;
      end
    end
    if (_T_3190) begin
      if (_T_2080) begin
        dat_out_bypass_data_11 <= dat_rsp_img_11;
      end else begin
        dat_out_bypass_data_11 <= dat_rsp_conv_11;
      end
    end
    if (_T_3191) begin
      if (_T_2080) begin
        dat_out_bypass_data_12 <= dat_rsp_img_12;
      end else begin
        dat_out_bypass_data_12 <= dat_rsp_conv_12;
      end
    end
    if (_T_3192) begin
      if (_T_2080) begin
        dat_out_bypass_data_13 <= dat_rsp_img_13;
      end else begin
        dat_out_bypass_data_13 <= dat_rsp_conv_13;
      end
    end
    if (_T_3193) begin
      if (_T_2080) begin
        dat_out_bypass_data_14 <= dat_rsp_img_14;
      end else begin
        dat_out_bypass_data_14 <= dat_rsp_conv_14;
      end
    end
    if (_T_3194) begin
      if (_T_2080) begin
        dat_out_bypass_data_15 <= dat_rsp_img_15;
      end else begin
        dat_out_bypass_data_15 <= dat_rsp_conv_15;
      end
    end
    if (_T_3195) begin
      if (_T_2080) begin
        dat_out_bypass_data_16 <= dat_rsp_img_16;
      end else begin
        dat_out_bypass_data_16 <= dat_rsp_conv_16;
      end
    end
    if (_T_3196) begin
      if (_T_2080) begin
        dat_out_bypass_data_17 <= dat_rsp_img_17;
      end else begin
        dat_out_bypass_data_17 <= dat_rsp_conv_17;
      end
    end
    if (_T_3197) begin
      if (_T_2080) begin
        dat_out_bypass_data_18 <= dat_rsp_img_18;
      end else begin
        dat_out_bypass_data_18 <= dat_rsp_conv_18;
      end
    end
    if (_T_3198) begin
      if (_T_2080) begin
        dat_out_bypass_data_19 <= dat_rsp_img_19;
      end else begin
        dat_out_bypass_data_19 <= dat_rsp_conv_19;
      end
    end
    if (_T_3199) begin
      if (_T_2080) begin
        dat_out_bypass_data_20 <= dat_rsp_img_20;
      end else begin
        dat_out_bypass_data_20 <= dat_rsp_conv_20;
      end
    end
    if (_T_3200) begin
      if (_T_2080) begin
        dat_out_bypass_data_21 <= dat_rsp_img_21;
      end else begin
        dat_out_bypass_data_21 <= dat_rsp_conv_21;
      end
    end
    if (_T_3201) begin
      if (_T_2080) begin
        dat_out_bypass_data_22 <= dat_rsp_img_22;
      end else begin
        dat_out_bypass_data_22 <= dat_rsp_conv_22;
      end
    end
    if (_T_3202) begin
      if (_T_2080) begin
        dat_out_bypass_data_23 <= dat_rsp_img_23;
      end else begin
        dat_out_bypass_data_23 <= dat_rsp_conv_23;
      end
    end
    if (_T_3203) begin
      if (_T_2080) begin
        dat_out_bypass_data_24 <= dat_rsp_img_24;
      end else begin
        dat_out_bypass_data_24 <= dat_rsp_conv_24;
      end
    end
    if (_T_3204) begin
      if (_T_2080) begin
        dat_out_bypass_data_25 <= dat_rsp_img_25;
      end else begin
        dat_out_bypass_data_25 <= dat_rsp_conv_25;
      end
    end
    if (_T_3205) begin
      if (_T_2080) begin
        dat_out_bypass_data_26 <= dat_rsp_img_26;
      end else begin
        dat_out_bypass_data_26 <= dat_rsp_conv_26;
      end
    end
    if (_T_3206) begin
      if (_T_2080) begin
        dat_out_bypass_data_27 <= dat_rsp_img_27;
      end else begin
        dat_out_bypass_data_27 <= dat_rsp_conv_27;
      end
    end
    if (_T_3207) begin
      if (_T_2080) begin
        dat_out_bypass_data_28 <= dat_rsp_img_28;
      end else begin
        dat_out_bypass_data_28 <= dat_rsp_conv_28;
      end
    end
    if (_T_3208) begin
      if (_T_2080) begin
        dat_out_bypass_data_29 <= dat_rsp_img_29;
      end else begin
        dat_out_bypass_data_29 <= dat_rsp_conv_29;
      end
    end
    if (_T_3209) begin
      if (_T_2080) begin
        dat_out_bypass_data_30 <= dat_rsp_img_30;
      end else begin
        dat_out_bypass_data_30 <= dat_rsp_conv_30;
      end
    end
    if (_T_3210) begin
      if (_T_2080) begin
        dat_out_bypass_data_31 <= dat_rsp_img_31;
      end else begin
        dat_out_bypass_data_31 <= dat_rsp_conv_31;
      end
    end
    if (_T_3211) begin
      if (_T_2080) begin
        dat_out_bypass_data_32 <= dat_rsp_img_32;
      end else begin
        dat_out_bypass_data_32 <= dat_rsp_conv_32;
      end
    end
    if (_T_3212) begin
      if (_T_2080) begin
        dat_out_bypass_data_33 <= dat_rsp_img_33;
      end else begin
        dat_out_bypass_data_33 <= dat_rsp_conv_33;
      end
    end
    if (_T_3213) begin
      if (_T_2080) begin
        dat_out_bypass_data_34 <= dat_rsp_img_34;
      end else begin
        dat_out_bypass_data_34 <= dat_rsp_conv_34;
      end
    end
    if (_T_3214) begin
      if (_T_2080) begin
        dat_out_bypass_data_35 <= dat_rsp_img_35;
      end else begin
        dat_out_bypass_data_35 <= dat_rsp_conv_35;
      end
    end
    if (_T_3215) begin
      if (_T_2080) begin
        dat_out_bypass_data_36 <= dat_rsp_img_36;
      end else begin
        dat_out_bypass_data_36 <= dat_rsp_conv_36;
      end
    end
    if (_T_3216) begin
      if (_T_2080) begin
        dat_out_bypass_data_37 <= dat_rsp_img_37;
      end else begin
        dat_out_bypass_data_37 <= dat_rsp_conv_37;
      end
    end
    if (_T_3217) begin
      if (_T_2080) begin
        dat_out_bypass_data_38 <= dat_rsp_img_38;
      end else begin
        dat_out_bypass_data_38 <= dat_rsp_conv_38;
      end
    end
    if (_T_3218) begin
      if (_T_2080) begin
        dat_out_bypass_data_39 <= dat_rsp_img_39;
      end else begin
        dat_out_bypass_data_39 <= dat_rsp_conv_39;
      end
    end
    if (_T_3219) begin
      if (_T_2080) begin
        dat_out_bypass_data_40 <= dat_rsp_img_40;
      end else begin
        dat_out_bypass_data_40 <= dat_rsp_conv_40;
      end
    end
    if (_T_3220) begin
      if (_T_2080) begin
        dat_out_bypass_data_41 <= dat_rsp_img_41;
      end else begin
        dat_out_bypass_data_41 <= dat_rsp_conv_41;
      end
    end
    if (_T_3221) begin
      if (_T_2080) begin
        dat_out_bypass_data_42 <= dat_rsp_img_42;
      end else begin
        dat_out_bypass_data_42 <= dat_rsp_conv_42;
      end
    end
    if (_T_3222) begin
      if (_T_2080) begin
        dat_out_bypass_data_43 <= dat_rsp_img_43;
      end else begin
        dat_out_bypass_data_43 <= dat_rsp_conv_43;
      end
    end
    if (_T_3223) begin
      if (_T_2080) begin
        dat_out_bypass_data_44 <= dat_rsp_img_44;
      end else begin
        dat_out_bypass_data_44 <= dat_rsp_conv_44;
      end
    end
    if (_T_3224) begin
      if (_T_2080) begin
        dat_out_bypass_data_45 <= dat_rsp_img_45;
      end else begin
        dat_out_bypass_data_45 <= dat_rsp_conv_45;
      end
    end
    if (_T_3225) begin
      if (_T_2080) begin
        dat_out_bypass_data_46 <= dat_rsp_img_46;
      end else begin
        dat_out_bypass_data_46 <= dat_rsp_conv_46;
      end
    end
    if (_T_3226) begin
      if (_T_2080) begin
        dat_out_bypass_data_47 <= dat_rsp_img_47;
      end else begin
        dat_out_bypass_data_47 <= dat_rsp_conv_47;
      end
    end
    if (_T_3227) begin
      if (_T_2080) begin
        dat_out_bypass_data_48 <= dat_rsp_img_48;
      end else begin
        dat_out_bypass_data_48 <= dat_rsp_conv_48;
      end
    end
    if (_T_3228) begin
      if (_T_2080) begin
        dat_out_bypass_data_49 <= dat_rsp_img_49;
      end else begin
        dat_out_bypass_data_49 <= dat_rsp_conv_49;
      end
    end
    if (_T_3229) begin
      if (_T_2080) begin
        dat_out_bypass_data_50 <= dat_rsp_img_50;
      end else begin
        dat_out_bypass_data_50 <= dat_rsp_conv_50;
      end
    end
    if (_T_3230) begin
      if (_T_2080) begin
        dat_out_bypass_data_51 <= dat_rsp_img_51;
      end else begin
        dat_out_bypass_data_51 <= dat_rsp_conv_51;
      end
    end
    if (_T_3231) begin
      if (_T_2080) begin
        dat_out_bypass_data_52 <= dat_rsp_img_52;
      end else begin
        dat_out_bypass_data_52 <= dat_rsp_conv_52;
      end
    end
    if (_T_3232) begin
      if (_T_2080) begin
        dat_out_bypass_data_53 <= dat_rsp_img_53;
      end else begin
        dat_out_bypass_data_53 <= dat_rsp_conv_53;
      end
    end
    if (_T_3233) begin
      if (_T_2080) begin
        dat_out_bypass_data_54 <= dat_rsp_img_54;
      end else begin
        dat_out_bypass_data_54 <= dat_rsp_conv_54;
      end
    end
    if (_T_3234) begin
      if (_T_2080) begin
        dat_out_bypass_data_55 <= dat_rsp_img_55;
      end else begin
        dat_out_bypass_data_55 <= dat_rsp_conv_55;
      end
    end
    if (_T_3235) begin
      if (_T_2080) begin
        dat_out_bypass_data_56 <= dat_rsp_img_56;
      end else begin
        dat_out_bypass_data_56 <= dat_rsp_conv_56;
      end
    end
    if (_T_3236) begin
      if (_T_2080) begin
        dat_out_bypass_data_57 <= dat_rsp_img_57;
      end else begin
        dat_out_bypass_data_57 <= dat_rsp_conv_57;
      end
    end
    if (_T_3237) begin
      if (_T_2080) begin
        dat_out_bypass_data_58 <= dat_rsp_img_58;
      end else begin
        dat_out_bypass_data_58 <= dat_rsp_conv_58;
      end
    end
    if (_T_3238) begin
      if (_T_2080) begin
        dat_out_bypass_data_59 <= dat_rsp_img_59;
      end else begin
        dat_out_bypass_data_59 <= dat_rsp_conv_59;
      end
    end
    if (_T_3239) begin
      if (_T_2080) begin
        dat_out_bypass_data_60 <= dat_rsp_img_60;
      end else begin
        dat_out_bypass_data_60 <= dat_rsp_conv_60;
      end
    end
    if (_T_3240) begin
      if (_T_2080) begin
        dat_out_bypass_data_61 <= dat_rsp_img_61;
      end else begin
        dat_out_bypass_data_61 <= dat_rsp_conv_61;
      end
    end
    if (_T_3241) begin
      if (_T_2080) begin
        dat_out_bypass_data_62 <= dat_rsp_img_62;
      end else begin
        dat_out_bypass_data_62 <= dat_rsp_conv_62;
      end
    end
    if (_T_3242) begin
      if (_T_2080) begin
        dat_out_bypass_data_63 <= dat_rsp_img_63;
      end else begin
        dat_out_bypass_data_63 <= dat_rsp_conv_63;
      end
    end
    if (_T_207) begin
      _T_3147 <= 1'h0;
    end else begin
      _T_3147 <= dat_rsp_pvld;
    end
    if (_T_207) begin
      _T_3150 <= 1'h0;
    end else begin
      _T_3150 <= _T_3147;
    end
    if (_T_207) begin
      _T_3153 <= 1'h0;
    end else begin
      _T_3153 <= _T_3150;
    end
    if (_T_207) begin
      _T_3156 <= 1'h0;
    end else begin
      _T_3156 <= _T_3153;
    end
    if (_T_207) begin
      _T_3159 <= 1'h0;
    end else begin
      _T_3159 <= _T_3156;
    end
    if (_T_207) begin
      _T_3164 <= 9'h0;
    end else begin
      if (dat_rsp_pvld) begin
        _T_3164 <= dat_rsp_flag;
      end
    end
    if (_T_207) begin
      _T_3167 <= 9'h0;
    end else begin
      if (_T_3147) begin
        _T_3167 <= _T_3164;
      end
    end
    if (_T_207) begin
      _T_3170 <= 9'h0;
    end else begin
      if (_T_3150) begin
        _T_3170 <= _T_3167;
      end
    end
    if (_T_207) begin
      _T_3173 <= 9'h0;
    end else begin
      if (_T_3153) begin
        _T_3173 <= _T_3170;
      end
    end
    if (_T_207) begin
      _T_3176 <= 9'h0;
    end else begin
      if (_T_3156) begin
        _T_3176 <= _T_3173;
      end
    end
    if (_T_207) begin
      dl_out_pvld <= 1'h0;
    end else begin
      dl_out_pvld <= dat_out_pvld;
    end
    if (_T_207) begin
      dl_out_mask_0 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_0 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_0 <= 1'h0;
          end else begin
            dl_out_mask_0 <= dat_out_bypass_mask_0;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_1 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_1 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_1 <= 1'h0;
          end else begin
            dl_out_mask_1 <= dat_out_bypass_mask_1;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_2 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_2 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_2 <= 1'h0;
          end else begin
            dl_out_mask_2 <= dat_out_bypass_mask_2;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_3 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_3 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_3 <= 1'h0;
          end else begin
            dl_out_mask_3 <= dat_out_bypass_mask_3;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_4 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_4 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_4 <= 1'h0;
          end else begin
            dl_out_mask_4 <= dat_out_bypass_mask_4;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_5 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_5 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_5 <= 1'h0;
          end else begin
            dl_out_mask_5 <= dat_out_bypass_mask_5;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_6 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_6 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_6 <= 1'h0;
          end else begin
            dl_out_mask_6 <= dat_out_bypass_mask_6;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_7 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_7 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_7 <= 1'h0;
          end else begin
            dl_out_mask_7 <= dat_out_bypass_mask_7;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_8 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_8 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_8 <= 1'h0;
          end else begin
            dl_out_mask_8 <= dat_out_bypass_mask_8;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_9 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_9 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_9 <= 1'h0;
          end else begin
            dl_out_mask_9 <= dat_out_bypass_mask_9;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_10 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_10 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_10 <= 1'h0;
          end else begin
            dl_out_mask_10 <= dat_out_bypass_mask_10;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_11 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_11 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_11 <= 1'h0;
          end else begin
            dl_out_mask_11 <= dat_out_bypass_mask_11;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_12 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_12 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_12 <= 1'h0;
          end else begin
            dl_out_mask_12 <= dat_out_bypass_mask_12;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_13 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_13 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_13 <= 1'h0;
          end else begin
            dl_out_mask_13 <= dat_out_bypass_mask_13;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_14 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_14 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_14 <= 1'h0;
          end else begin
            dl_out_mask_14 <= dat_out_bypass_mask_14;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_15 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_15 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_15 <= 1'h0;
          end else begin
            dl_out_mask_15 <= dat_out_bypass_mask_15;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_16 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_16 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_16 <= 1'h0;
          end else begin
            dl_out_mask_16 <= dat_out_bypass_mask_16;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_17 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_17 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_17 <= 1'h0;
          end else begin
            dl_out_mask_17 <= dat_out_bypass_mask_17;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_18 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_18 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_18 <= 1'h0;
          end else begin
            dl_out_mask_18 <= dat_out_bypass_mask_18;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_19 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_19 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_19 <= 1'h0;
          end else begin
            dl_out_mask_19 <= dat_out_bypass_mask_19;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_20 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_20 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_20 <= 1'h0;
          end else begin
            dl_out_mask_20 <= dat_out_bypass_mask_20;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_21 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_21 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_21 <= 1'h0;
          end else begin
            dl_out_mask_21 <= dat_out_bypass_mask_21;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_22 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_22 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_22 <= 1'h0;
          end else begin
            dl_out_mask_22 <= dat_out_bypass_mask_22;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_23 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_23 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_23 <= 1'h0;
          end else begin
            dl_out_mask_23 <= dat_out_bypass_mask_23;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_24 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_24 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_24 <= 1'h0;
          end else begin
            dl_out_mask_24 <= dat_out_bypass_mask_24;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_25 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_25 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_25 <= 1'h0;
          end else begin
            dl_out_mask_25 <= dat_out_bypass_mask_25;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_26 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_26 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_26 <= 1'h0;
          end else begin
            dl_out_mask_26 <= dat_out_bypass_mask_26;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_27 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_27 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_27 <= 1'h0;
          end else begin
            dl_out_mask_27 <= dat_out_bypass_mask_27;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_28 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_28 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_28 <= 1'h0;
          end else begin
            dl_out_mask_28 <= dat_out_bypass_mask_28;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_29 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_29 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_29 <= 1'h0;
          end else begin
            dl_out_mask_29 <= dat_out_bypass_mask_29;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_30 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_30 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_30 <= 1'h0;
          end else begin
            dl_out_mask_30 <= dat_out_bypass_mask_30;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_31 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_31 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_31 <= 1'h0;
          end else begin
            dl_out_mask_31 <= dat_out_bypass_mask_31;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_32 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_32 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_32 <= 1'h0;
          end else begin
            dl_out_mask_32 <= dat_out_bypass_mask_32;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_33 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_33 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_33 <= 1'h0;
          end else begin
            dl_out_mask_33 <= dat_out_bypass_mask_33;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_34 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_34 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_34 <= 1'h0;
          end else begin
            dl_out_mask_34 <= dat_out_bypass_mask_34;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_35 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_35 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_35 <= 1'h0;
          end else begin
            dl_out_mask_35 <= dat_out_bypass_mask_35;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_36 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_36 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_36 <= 1'h0;
          end else begin
            dl_out_mask_36 <= dat_out_bypass_mask_36;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_37 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_37 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_37 <= 1'h0;
          end else begin
            dl_out_mask_37 <= dat_out_bypass_mask_37;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_38 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_38 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_38 <= 1'h0;
          end else begin
            dl_out_mask_38 <= dat_out_bypass_mask_38;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_39 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_39 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_39 <= 1'h0;
          end else begin
            dl_out_mask_39 <= dat_out_bypass_mask_39;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_40 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_40 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_40 <= 1'h0;
          end else begin
            dl_out_mask_40 <= dat_out_bypass_mask_40;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_41 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_41 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_41 <= 1'h0;
          end else begin
            dl_out_mask_41 <= dat_out_bypass_mask_41;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_42 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_42 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_42 <= 1'h0;
          end else begin
            dl_out_mask_42 <= dat_out_bypass_mask_42;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_43 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_43 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_43 <= 1'h0;
          end else begin
            dl_out_mask_43 <= dat_out_bypass_mask_43;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_44 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_44 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_44 <= 1'h0;
          end else begin
            dl_out_mask_44 <= dat_out_bypass_mask_44;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_45 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_45 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_45 <= 1'h0;
          end else begin
            dl_out_mask_45 <= dat_out_bypass_mask_45;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_46 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_46 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_46 <= 1'h0;
          end else begin
            dl_out_mask_46 <= dat_out_bypass_mask_46;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_47 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_47 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_47 <= 1'h0;
          end else begin
            dl_out_mask_47 <= dat_out_bypass_mask_47;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_48 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_48 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_48 <= 1'h0;
          end else begin
            dl_out_mask_48 <= dat_out_bypass_mask_48;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_49 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_49 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_49 <= 1'h0;
          end else begin
            dl_out_mask_49 <= dat_out_bypass_mask_49;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_50 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_50 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_50 <= 1'h0;
          end else begin
            dl_out_mask_50 <= dat_out_bypass_mask_50;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_51 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_51 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_51 <= 1'h0;
          end else begin
            dl_out_mask_51 <= dat_out_bypass_mask_51;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_52 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_52 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_52 <= 1'h0;
          end else begin
            dl_out_mask_52 <= dat_out_bypass_mask_52;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_53 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_53 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_53 <= 1'h0;
          end else begin
            dl_out_mask_53 <= dat_out_bypass_mask_53;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_54 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_54 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_54 <= 1'h0;
          end else begin
            dl_out_mask_54 <= dat_out_bypass_mask_54;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_55 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_55 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_55 <= 1'h0;
          end else begin
            dl_out_mask_55 <= dat_out_bypass_mask_55;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_56 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_56 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_56 <= 1'h0;
          end else begin
            dl_out_mask_56 <= dat_out_bypass_mask_56;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_57 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_57 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_57 <= 1'h0;
          end else begin
            dl_out_mask_57 <= dat_out_bypass_mask_57;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_58 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_58 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_58 <= 1'h0;
          end else begin
            dl_out_mask_58 <= dat_out_bypass_mask_58;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_59 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_59 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_59 <= 1'h0;
          end else begin
            dl_out_mask_59 <= dat_out_bypass_mask_59;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_60 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_60 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_60 <= 1'h0;
          end else begin
            dl_out_mask_60 <= dat_out_bypass_mask_60;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_61 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_61 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_61 <= 1'h0;
          end else begin
            dl_out_mask_61 <= dat_out_bypass_mask_61;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_62 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_62 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_62 <= 1'h0;
          end else begin
            dl_out_mask_62 <= dat_out_bypass_mask_62;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_mask_63 <= 1'h0;
    end else begin
      if (_T_4575) begin
        if (_T_4176) begin
          dl_out_mask_63 <= 1'h0;
        end else begin
          if (_T_4311) begin
            dl_out_mask_63 <= 1'h0;
          end else begin
            dl_out_mask_63 <= dat_out_bypass_mask_63;
          end
        end
      end
    end
    if (_T_207) begin
      dl_out_flag <= 9'h0;
    end else begin
      if (dat_out_pvld) begin
        dl_out_flag <= dat_out_flag;
      end
    end
    if (dat_out_mask_0) begin
      if (_T_4044) begin
        dl_out_data_0 <= 8'h0;
      end else begin
        dl_out_data_0 <= dat_out_bypass_data_0;
      end
    end
    if (dat_out_mask_1) begin
      if (_T_4044) begin
        dl_out_data_1 <= 8'h0;
      end else begin
        dl_out_data_1 <= dat_out_bypass_data_1;
      end
    end
    if (dat_out_mask_2) begin
      if (_T_4044) begin
        dl_out_data_2 <= 8'h0;
      end else begin
        dl_out_data_2 <= dat_out_bypass_data_2;
      end
    end
    if (dat_out_mask_3) begin
      if (_T_4044) begin
        dl_out_data_3 <= 8'h0;
      end else begin
        dl_out_data_3 <= dat_out_bypass_data_3;
      end
    end
    if (dat_out_mask_4) begin
      if (_T_4044) begin
        dl_out_data_4 <= 8'h0;
      end else begin
        dl_out_data_4 <= dat_out_bypass_data_4;
      end
    end
    if (dat_out_mask_5) begin
      if (_T_4044) begin
        dl_out_data_5 <= 8'h0;
      end else begin
        dl_out_data_5 <= dat_out_bypass_data_5;
      end
    end
    if (dat_out_mask_6) begin
      if (_T_4044) begin
        dl_out_data_6 <= 8'h0;
      end else begin
        dl_out_data_6 <= dat_out_bypass_data_6;
      end
    end
    if (dat_out_mask_7) begin
      if (_T_4044) begin
        dl_out_data_7 <= 8'h0;
      end else begin
        dl_out_data_7 <= dat_out_bypass_data_7;
      end
    end
    if (dat_out_mask_8) begin
      if (_T_4044) begin
        dl_out_data_8 <= 8'h0;
      end else begin
        dl_out_data_8 <= dat_out_bypass_data_8;
      end
    end
    if (dat_out_mask_9) begin
      if (_T_4044) begin
        dl_out_data_9 <= 8'h0;
      end else begin
        dl_out_data_9 <= dat_out_bypass_data_9;
      end
    end
    if (dat_out_mask_10) begin
      if (_T_4044) begin
        dl_out_data_10 <= 8'h0;
      end else begin
        dl_out_data_10 <= dat_out_bypass_data_10;
      end
    end
    if (dat_out_mask_11) begin
      if (_T_4044) begin
        dl_out_data_11 <= 8'h0;
      end else begin
        dl_out_data_11 <= dat_out_bypass_data_11;
      end
    end
    if (dat_out_mask_12) begin
      if (_T_4044) begin
        dl_out_data_12 <= 8'h0;
      end else begin
        dl_out_data_12 <= dat_out_bypass_data_12;
      end
    end
    if (dat_out_mask_13) begin
      if (_T_4044) begin
        dl_out_data_13 <= 8'h0;
      end else begin
        dl_out_data_13 <= dat_out_bypass_data_13;
      end
    end
    if (dat_out_mask_14) begin
      if (_T_4044) begin
        dl_out_data_14 <= 8'h0;
      end else begin
        dl_out_data_14 <= dat_out_bypass_data_14;
      end
    end
    if (dat_out_mask_15) begin
      if (_T_4044) begin
        dl_out_data_15 <= 8'h0;
      end else begin
        dl_out_data_15 <= dat_out_bypass_data_15;
      end
    end
    if (dat_out_mask_16) begin
      if (_T_4044) begin
        dl_out_data_16 <= 8'h0;
      end else begin
        dl_out_data_16 <= dat_out_bypass_data_16;
      end
    end
    if (dat_out_mask_17) begin
      if (_T_4044) begin
        dl_out_data_17 <= 8'h0;
      end else begin
        dl_out_data_17 <= dat_out_bypass_data_17;
      end
    end
    if (dat_out_mask_18) begin
      if (_T_4044) begin
        dl_out_data_18 <= 8'h0;
      end else begin
        dl_out_data_18 <= dat_out_bypass_data_18;
      end
    end
    if (dat_out_mask_19) begin
      if (_T_4044) begin
        dl_out_data_19 <= 8'h0;
      end else begin
        dl_out_data_19 <= dat_out_bypass_data_19;
      end
    end
    if (dat_out_mask_20) begin
      if (_T_4044) begin
        dl_out_data_20 <= 8'h0;
      end else begin
        dl_out_data_20 <= dat_out_bypass_data_20;
      end
    end
    if (dat_out_mask_21) begin
      if (_T_4044) begin
        dl_out_data_21 <= 8'h0;
      end else begin
        dl_out_data_21 <= dat_out_bypass_data_21;
      end
    end
    if (dat_out_mask_22) begin
      if (_T_4044) begin
        dl_out_data_22 <= 8'h0;
      end else begin
        dl_out_data_22 <= dat_out_bypass_data_22;
      end
    end
    if (dat_out_mask_23) begin
      if (_T_4044) begin
        dl_out_data_23 <= 8'h0;
      end else begin
        dl_out_data_23 <= dat_out_bypass_data_23;
      end
    end
    if (dat_out_mask_24) begin
      if (_T_4044) begin
        dl_out_data_24 <= 8'h0;
      end else begin
        dl_out_data_24 <= dat_out_bypass_data_24;
      end
    end
    if (dat_out_mask_25) begin
      if (_T_4044) begin
        dl_out_data_25 <= 8'h0;
      end else begin
        dl_out_data_25 <= dat_out_bypass_data_25;
      end
    end
    if (dat_out_mask_26) begin
      if (_T_4044) begin
        dl_out_data_26 <= 8'h0;
      end else begin
        dl_out_data_26 <= dat_out_bypass_data_26;
      end
    end
    if (dat_out_mask_27) begin
      if (_T_4044) begin
        dl_out_data_27 <= 8'h0;
      end else begin
        dl_out_data_27 <= dat_out_bypass_data_27;
      end
    end
    if (dat_out_mask_28) begin
      if (_T_4044) begin
        dl_out_data_28 <= 8'h0;
      end else begin
        dl_out_data_28 <= dat_out_bypass_data_28;
      end
    end
    if (dat_out_mask_29) begin
      if (_T_4044) begin
        dl_out_data_29 <= 8'h0;
      end else begin
        dl_out_data_29 <= dat_out_bypass_data_29;
      end
    end
    if (dat_out_mask_30) begin
      if (_T_4044) begin
        dl_out_data_30 <= 8'h0;
      end else begin
        dl_out_data_30 <= dat_out_bypass_data_30;
      end
    end
    if (dat_out_mask_31) begin
      if (_T_4044) begin
        dl_out_data_31 <= 8'h0;
      end else begin
        dl_out_data_31 <= dat_out_bypass_data_31;
      end
    end
    if (dat_out_mask_32) begin
      if (_T_4044) begin
        dl_out_data_32 <= 8'h0;
      end else begin
        dl_out_data_32 <= dat_out_bypass_data_32;
      end
    end
    if (dat_out_mask_33) begin
      if (_T_4044) begin
        dl_out_data_33 <= 8'h0;
      end else begin
        dl_out_data_33 <= dat_out_bypass_data_33;
      end
    end
    if (dat_out_mask_34) begin
      if (_T_4044) begin
        dl_out_data_34 <= 8'h0;
      end else begin
        dl_out_data_34 <= dat_out_bypass_data_34;
      end
    end
    if (dat_out_mask_35) begin
      if (_T_4044) begin
        dl_out_data_35 <= 8'h0;
      end else begin
        dl_out_data_35 <= dat_out_bypass_data_35;
      end
    end
    if (dat_out_mask_36) begin
      if (_T_4044) begin
        dl_out_data_36 <= 8'h0;
      end else begin
        dl_out_data_36 <= dat_out_bypass_data_36;
      end
    end
    if (dat_out_mask_37) begin
      if (_T_4044) begin
        dl_out_data_37 <= 8'h0;
      end else begin
        dl_out_data_37 <= dat_out_bypass_data_37;
      end
    end
    if (dat_out_mask_38) begin
      if (_T_4044) begin
        dl_out_data_38 <= 8'h0;
      end else begin
        dl_out_data_38 <= dat_out_bypass_data_38;
      end
    end
    if (dat_out_mask_39) begin
      if (_T_4044) begin
        dl_out_data_39 <= 8'h0;
      end else begin
        dl_out_data_39 <= dat_out_bypass_data_39;
      end
    end
    if (dat_out_mask_40) begin
      if (_T_4044) begin
        dl_out_data_40 <= 8'h0;
      end else begin
        dl_out_data_40 <= dat_out_bypass_data_40;
      end
    end
    if (dat_out_mask_41) begin
      if (_T_4044) begin
        dl_out_data_41 <= 8'h0;
      end else begin
        dl_out_data_41 <= dat_out_bypass_data_41;
      end
    end
    if (dat_out_mask_42) begin
      if (_T_4044) begin
        dl_out_data_42 <= 8'h0;
      end else begin
        dl_out_data_42 <= dat_out_bypass_data_42;
      end
    end
    if (dat_out_mask_43) begin
      if (_T_4044) begin
        dl_out_data_43 <= 8'h0;
      end else begin
        dl_out_data_43 <= dat_out_bypass_data_43;
      end
    end
    if (dat_out_mask_44) begin
      if (_T_4044) begin
        dl_out_data_44 <= 8'h0;
      end else begin
        dl_out_data_44 <= dat_out_bypass_data_44;
      end
    end
    if (dat_out_mask_45) begin
      if (_T_4044) begin
        dl_out_data_45 <= 8'h0;
      end else begin
        dl_out_data_45 <= dat_out_bypass_data_45;
      end
    end
    if (dat_out_mask_46) begin
      if (_T_4044) begin
        dl_out_data_46 <= 8'h0;
      end else begin
        dl_out_data_46 <= dat_out_bypass_data_46;
      end
    end
    if (dat_out_mask_47) begin
      if (_T_4044) begin
        dl_out_data_47 <= 8'h0;
      end else begin
        dl_out_data_47 <= dat_out_bypass_data_47;
      end
    end
    if (dat_out_mask_48) begin
      if (_T_4044) begin
        dl_out_data_48 <= 8'h0;
      end else begin
        dl_out_data_48 <= dat_out_bypass_data_48;
      end
    end
    if (dat_out_mask_49) begin
      if (_T_4044) begin
        dl_out_data_49 <= 8'h0;
      end else begin
        dl_out_data_49 <= dat_out_bypass_data_49;
      end
    end
    if (dat_out_mask_50) begin
      if (_T_4044) begin
        dl_out_data_50 <= 8'h0;
      end else begin
        dl_out_data_50 <= dat_out_bypass_data_50;
      end
    end
    if (dat_out_mask_51) begin
      if (_T_4044) begin
        dl_out_data_51 <= 8'h0;
      end else begin
        dl_out_data_51 <= dat_out_bypass_data_51;
      end
    end
    if (dat_out_mask_52) begin
      if (_T_4044) begin
        dl_out_data_52 <= 8'h0;
      end else begin
        dl_out_data_52 <= dat_out_bypass_data_52;
      end
    end
    if (dat_out_mask_53) begin
      if (_T_4044) begin
        dl_out_data_53 <= 8'h0;
      end else begin
        dl_out_data_53 <= dat_out_bypass_data_53;
      end
    end
    if (dat_out_mask_54) begin
      if (_T_4044) begin
        dl_out_data_54 <= 8'h0;
      end else begin
        dl_out_data_54 <= dat_out_bypass_data_54;
      end
    end
    if (dat_out_mask_55) begin
      if (_T_4044) begin
        dl_out_data_55 <= 8'h0;
      end else begin
        dl_out_data_55 <= dat_out_bypass_data_55;
      end
    end
    if (dat_out_mask_56) begin
      if (_T_4044) begin
        dl_out_data_56 <= 8'h0;
      end else begin
        dl_out_data_56 <= dat_out_bypass_data_56;
      end
    end
    if (dat_out_mask_57) begin
      if (_T_4044) begin
        dl_out_data_57 <= 8'h0;
      end else begin
        dl_out_data_57 <= dat_out_bypass_data_57;
      end
    end
    if (dat_out_mask_58) begin
      if (_T_4044) begin
        dl_out_data_58 <= 8'h0;
      end else begin
        dl_out_data_58 <= dat_out_bypass_data_58;
      end
    end
    if (dat_out_mask_59) begin
      if (_T_4044) begin
        dl_out_data_59 <= 8'h0;
      end else begin
        dl_out_data_59 <= dat_out_bypass_data_59;
      end
    end
    if (dat_out_mask_60) begin
      if (_T_4044) begin
        dl_out_data_60 <= 8'h0;
      end else begin
        dl_out_data_60 <= dat_out_bypass_data_60;
      end
    end
    if (dat_out_mask_61) begin
      if (_T_4044) begin
        dl_out_data_61 <= 8'h0;
      end else begin
        dl_out_data_61 <= dat_out_bypass_data_61;
      end
    end
    if (dat_out_mask_62) begin
      if (_T_4044) begin
        dl_out_data_62 <= 8'h0;
      end else begin
        dl_out_data_62 <= dat_out_bypass_data_62;
      end
    end
    if (dat_out_mask_63) begin
      if (_T_4044) begin
        dl_out_data_63 <= 8'h0;
      end else begin
        dl_out_data_63 <= dat_out_bypass_data_63;
      end
    end
    if (_T_207) begin
      dl_out_pvld_d1 <= 1'h0;
    end else begin
      dl_out_pvld_d1 <= dl_out_pvld;
    end
    if (_T_207) begin
      _T_4582 <= 1'h0;
    end else begin
      _T_4582 <= dl_out_pvld;
    end
    if (_T_207) begin
      _T_4585 <= 1'h0;
    end else begin
      _T_4585 <= dl_out_pvld;
    end
    if (_T_207) begin
      _T_4589 <= 9'h0;
    end else begin
      if (_T_4587) begin
        if (_T_4578) begin
          _T_4589 <= 9'h0;
        end else begin
          _T_4589 <= dl_out_flag;
        end
      end
    end
    if (_T_207) begin
      _T_4593 <= 9'h0;
    end else begin
      if (_T_4587) begin
        if (_T_4578) begin
          _T_4593 <= 9'h0;
        end else begin
          _T_4593 <= dl_out_flag;
        end
      end
    end
    if (_T_207) begin
      _T_4861_0 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_0 <= dl_out_mask_0;
      end
    end
    if (_T_207) begin
      _T_4861_1 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_1 <= dl_out_mask_1;
      end
    end
    if (_T_207) begin
      _T_4861_2 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_2 <= dl_out_mask_2;
      end
    end
    if (_T_207) begin
      _T_4861_3 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_3 <= dl_out_mask_3;
      end
    end
    if (_T_207) begin
      _T_4861_4 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_4 <= dl_out_mask_4;
      end
    end
    if (_T_207) begin
      _T_4861_5 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_5 <= dl_out_mask_5;
      end
    end
    if (_T_207) begin
      _T_4861_6 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_6 <= dl_out_mask_6;
      end
    end
    if (_T_207) begin
      _T_4861_7 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_7 <= dl_out_mask_7;
      end
    end
    if (_T_207) begin
      _T_4861_8 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_8 <= dl_out_mask_8;
      end
    end
    if (_T_207) begin
      _T_4861_9 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_9 <= dl_out_mask_9;
      end
    end
    if (_T_207) begin
      _T_4861_10 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_10 <= dl_out_mask_10;
      end
    end
    if (_T_207) begin
      _T_4861_11 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_11 <= dl_out_mask_11;
      end
    end
    if (_T_207) begin
      _T_4861_12 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_12 <= dl_out_mask_12;
      end
    end
    if (_T_207) begin
      _T_4861_13 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_13 <= dl_out_mask_13;
      end
    end
    if (_T_207) begin
      _T_4861_14 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_14 <= dl_out_mask_14;
      end
    end
    if (_T_207) begin
      _T_4861_15 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_15 <= dl_out_mask_15;
      end
    end
    if (_T_207) begin
      _T_4861_16 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_16 <= dl_out_mask_16;
      end
    end
    if (_T_207) begin
      _T_4861_17 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_17 <= dl_out_mask_17;
      end
    end
    if (_T_207) begin
      _T_4861_18 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_18 <= dl_out_mask_18;
      end
    end
    if (_T_207) begin
      _T_4861_19 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_19 <= dl_out_mask_19;
      end
    end
    if (_T_207) begin
      _T_4861_20 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_20 <= dl_out_mask_20;
      end
    end
    if (_T_207) begin
      _T_4861_21 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_21 <= dl_out_mask_21;
      end
    end
    if (_T_207) begin
      _T_4861_22 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_22 <= dl_out_mask_22;
      end
    end
    if (_T_207) begin
      _T_4861_23 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_23 <= dl_out_mask_23;
      end
    end
    if (_T_207) begin
      _T_4861_24 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_24 <= dl_out_mask_24;
      end
    end
    if (_T_207) begin
      _T_4861_25 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_25 <= dl_out_mask_25;
      end
    end
    if (_T_207) begin
      _T_4861_26 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_26 <= dl_out_mask_26;
      end
    end
    if (_T_207) begin
      _T_4861_27 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_27 <= dl_out_mask_27;
      end
    end
    if (_T_207) begin
      _T_4861_28 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_28 <= dl_out_mask_28;
      end
    end
    if (_T_207) begin
      _T_4861_29 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_29 <= dl_out_mask_29;
      end
    end
    if (_T_207) begin
      _T_4861_30 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_30 <= dl_out_mask_30;
      end
    end
    if (_T_207) begin
      _T_4861_31 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_31 <= dl_out_mask_31;
      end
    end
    if (_T_207) begin
      _T_4861_32 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_32 <= dl_out_mask_32;
      end
    end
    if (_T_207) begin
      _T_4861_33 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_33 <= dl_out_mask_33;
      end
    end
    if (_T_207) begin
      _T_4861_34 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_34 <= dl_out_mask_34;
      end
    end
    if (_T_207) begin
      _T_4861_35 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_35 <= dl_out_mask_35;
      end
    end
    if (_T_207) begin
      _T_4861_36 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_36 <= dl_out_mask_36;
      end
    end
    if (_T_207) begin
      _T_4861_37 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_37 <= dl_out_mask_37;
      end
    end
    if (_T_207) begin
      _T_4861_38 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_38 <= dl_out_mask_38;
      end
    end
    if (_T_207) begin
      _T_4861_39 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_39 <= dl_out_mask_39;
      end
    end
    if (_T_207) begin
      _T_4861_40 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_40 <= dl_out_mask_40;
      end
    end
    if (_T_207) begin
      _T_4861_41 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_41 <= dl_out_mask_41;
      end
    end
    if (_T_207) begin
      _T_4861_42 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_42 <= dl_out_mask_42;
      end
    end
    if (_T_207) begin
      _T_4861_43 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_43 <= dl_out_mask_43;
      end
    end
    if (_T_207) begin
      _T_4861_44 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_44 <= dl_out_mask_44;
      end
    end
    if (_T_207) begin
      _T_4861_45 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_45 <= dl_out_mask_45;
      end
    end
    if (_T_207) begin
      _T_4861_46 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_46 <= dl_out_mask_46;
      end
    end
    if (_T_207) begin
      _T_4861_47 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_47 <= dl_out_mask_47;
      end
    end
    if (_T_207) begin
      _T_4861_48 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_48 <= dl_out_mask_48;
      end
    end
    if (_T_207) begin
      _T_4861_49 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_49 <= dl_out_mask_49;
      end
    end
    if (_T_207) begin
      _T_4861_50 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_50 <= dl_out_mask_50;
      end
    end
    if (_T_207) begin
      _T_4861_51 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_51 <= dl_out_mask_51;
      end
    end
    if (_T_207) begin
      _T_4861_52 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_52 <= dl_out_mask_52;
      end
    end
    if (_T_207) begin
      _T_4861_53 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_53 <= dl_out_mask_53;
      end
    end
    if (_T_207) begin
      _T_4861_54 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_54 <= dl_out_mask_54;
      end
    end
    if (_T_207) begin
      _T_4861_55 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_55 <= dl_out_mask_55;
      end
    end
    if (_T_207) begin
      _T_4861_56 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_56 <= dl_out_mask_56;
      end
    end
    if (_T_207) begin
      _T_4861_57 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_57 <= dl_out_mask_57;
      end
    end
    if (_T_207) begin
      _T_4861_58 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_58 <= dl_out_mask_58;
      end
    end
    if (_T_207) begin
      _T_4861_59 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_59 <= dl_out_mask_59;
      end
    end
    if (_T_207) begin
      _T_4861_60 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_60 <= dl_out_mask_60;
      end
    end
    if (_T_207) begin
      _T_4861_61 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_61 <= dl_out_mask_61;
      end
    end
    if (_T_207) begin
      _T_4861_62 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_62 <= dl_out_mask_62;
      end
    end
    if (_T_207) begin
      _T_4861_63 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_4861_63 <= dl_out_mask_63;
      end
    end
    if (_T_207) begin
      _T_5388_0 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_0 <= dl_out_mask_0;
      end
    end
    if (_T_207) begin
      _T_5388_1 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_1 <= dl_out_mask_1;
      end
    end
    if (_T_207) begin
      _T_5388_2 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_2 <= dl_out_mask_2;
      end
    end
    if (_T_207) begin
      _T_5388_3 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_3 <= dl_out_mask_3;
      end
    end
    if (_T_207) begin
      _T_5388_4 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_4 <= dl_out_mask_4;
      end
    end
    if (_T_207) begin
      _T_5388_5 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_5 <= dl_out_mask_5;
      end
    end
    if (_T_207) begin
      _T_5388_6 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_6 <= dl_out_mask_6;
      end
    end
    if (_T_207) begin
      _T_5388_7 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_7 <= dl_out_mask_7;
      end
    end
    if (_T_207) begin
      _T_5388_8 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_8 <= dl_out_mask_8;
      end
    end
    if (_T_207) begin
      _T_5388_9 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_9 <= dl_out_mask_9;
      end
    end
    if (_T_207) begin
      _T_5388_10 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_10 <= dl_out_mask_10;
      end
    end
    if (_T_207) begin
      _T_5388_11 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_11 <= dl_out_mask_11;
      end
    end
    if (_T_207) begin
      _T_5388_12 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_12 <= dl_out_mask_12;
      end
    end
    if (_T_207) begin
      _T_5388_13 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_13 <= dl_out_mask_13;
      end
    end
    if (_T_207) begin
      _T_5388_14 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_14 <= dl_out_mask_14;
      end
    end
    if (_T_207) begin
      _T_5388_15 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_15 <= dl_out_mask_15;
      end
    end
    if (_T_207) begin
      _T_5388_16 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_16 <= dl_out_mask_16;
      end
    end
    if (_T_207) begin
      _T_5388_17 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_17 <= dl_out_mask_17;
      end
    end
    if (_T_207) begin
      _T_5388_18 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_18 <= dl_out_mask_18;
      end
    end
    if (_T_207) begin
      _T_5388_19 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_19 <= dl_out_mask_19;
      end
    end
    if (_T_207) begin
      _T_5388_20 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_20 <= dl_out_mask_20;
      end
    end
    if (_T_207) begin
      _T_5388_21 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_21 <= dl_out_mask_21;
      end
    end
    if (_T_207) begin
      _T_5388_22 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_22 <= dl_out_mask_22;
      end
    end
    if (_T_207) begin
      _T_5388_23 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_23 <= dl_out_mask_23;
      end
    end
    if (_T_207) begin
      _T_5388_24 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_24 <= dl_out_mask_24;
      end
    end
    if (_T_207) begin
      _T_5388_25 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_25 <= dl_out_mask_25;
      end
    end
    if (_T_207) begin
      _T_5388_26 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_26 <= dl_out_mask_26;
      end
    end
    if (_T_207) begin
      _T_5388_27 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_27 <= dl_out_mask_27;
      end
    end
    if (_T_207) begin
      _T_5388_28 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_28 <= dl_out_mask_28;
      end
    end
    if (_T_207) begin
      _T_5388_29 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_29 <= dl_out_mask_29;
      end
    end
    if (_T_207) begin
      _T_5388_30 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_30 <= dl_out_mask_30;
      end
    end
    if (_T_207) begin
      _T_5388_31 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_31 <= dl_out_mask_31;
      end
    end
    if (_T_207) begin
      _T_5388_32 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_32 <= dl_out_mask_32;
      end
    end
    if (_T_207) begin
      _T_5388_33 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_33 <= dl_out_mask_33;
      end
    end
    if (_T_207) begin
      _T_5388_34 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_34 <= dl_out_mask_34;
      end
    end
    if (_T_207) begin
      _T_5388_35 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_35 <= dl_out_mask_35;
      end
    end
    if (_T_207) begin
      _T_5388_36 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_36 <= dl_out_mask_36;
      end
    end
    if (_T_207) begin
      _T_5388_37 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_37 <= dl_out_mask_37;
      end
    end
    if (_T_207) begin
      _T_5388_38 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_38 <= dl_out_mask_38;
      end
    end
    if (_T_207) begin
      _T_5388_39 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_39 <= dl_out_mask_39;
      end
    end
    if (_T_207) begin
      _T_5388_40 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_40 <= dl_out_mask_40;
      end
    end
    if (_T_207) begin
      _T_5388_41 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_41 <= dl_out_mask_41;
      end
    end
    if (_T_207) begin
      _T_5388_42 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_42 <= dl_out_mask_42;
      end
    end
    if (_T_207) begin
      _T_5388_43 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_43 <= dl_out_mask_43;
      end
    end
    if (_T_207) begin
      _T_5388_44 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_44 <= dl_out_mask_44;
      end
    end
    if (_T_207) begin
      _T_5388_45 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_45 <= dl_out_mask_45;
      end
    end
    if (_T_207) begin
      _T_5388_46 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_46 <= dl_out_mask_46;
      end
    end
    if (_T_207) begin
      _T_5388_47 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_47 <= dl_out_mask_47;
      end
    end
    if (_T_207) begin
      _T_5388_48 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_48 <= dl_out_mask_48;
      end
    end
    if (_T_207) begin
      _T_5388_49 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_49 <= dl_out_mask_49;
      end
    end
    if (_T_207) begin
      _T_5388_50 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_50 <= dl_out_mask_50;
      end
    end
    if (_T_207) begin
      _T_5388_51 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_51 <= dl_out_mask_51;
      end
    end
    if (_T_207) begin
      _T_5388_52 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_52 <= dl_out_mask_52;
      end
    end
    if (_T_207) begin
      _T_5388_53 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_53 <= dl_out_mask_53;
      end
    end
    if (_T_207) begin
      _T_5388_54 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_54 <= dl_out_mask_54;
      end
    end
    if (_T_207) begin
      _T_5388_55 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_55 <= dl_out_mask_55;
      end
    end
    if (_T_207) begin
      _T_5388_56 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_56 <= dl_out_mask_56;
      end
    end
    if (_T_207) begin
      _T_5388_57 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_57 <= dl_out_mask_57;
      end
    end
    if (_T_207) begin
      _T_5388_58 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_58 <= dl_out_mask_58;
      end
    end
    if (_T_207) begin
      _T_5388_59 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_59 <= dl_out_mask_59;
      end
    end
    if (_T_207) begin
      _T_5388_60 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_60 <= dl_out_mask_60;
      end
    end
    if (_T_207) begin
      _T_5388_61 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_61 <= dl_out_mask_61;
      end
    end
    if (_T_207) begin
      _T_5388_62 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_62 <= dl_out_mask_62;
      end
    end
    if (_T_207) begin
      _T_5388_63 <= 1'h0;
    end else begin
      if (_T_4587) begin
        _T_5388_63 <= dl_out_mask_63;
      end
    end
    if (dl_out_mask_0) begin
      _T_5649 <= dl_out_data_0;
    end
    if (dl_out_mask_0) begin
      _T_5651 <= dl_out_data_0;
    end
    if (dl_out_mask_1) begin
      _T_5653 <= dl_out_data_1;
    end
    if (dl_out_mask_1) begin
      _T_5655 <= dl_out_data_1;
    end
    if (dl_out_mask_2) begin
      _T_5657 <= dl_out_data_2;
    end
    if (dl_out_mask_2) begin
      _T_5659 <= dl_out_data_2;
    end
    if (dl_out_mask_3) begin
      _T_5661 <= dl_out_data_3;
    end
    if (dl_out_mask_3) begin
      _T_5663 <= dl_out_data_3;
    end
    if (dl_out_mask_4) begin
      _T_5665 <= dl_out_data_4;
    end
    if (dl_out_mask_4) begin
      _T_5667 <= dl_out_data_4;
    end
    if (dl_out_mask_5) begin
      _T_5669 <= dl_out_data_5;
    end
    if (dl_out_mask_5) begin
      _T_5671 <= dl_out_data_5;
    end
    if (dl_out_mask_6) begin
      _T_5673 <= dl_out_data_6;
    end
    if (dl_out_mask_6) begin
      _T_5675 <= dl_out_data_6;
    end
    if (dl_out_mask_7) begin
      _T_5677 <= dl_out_data_7;
    end
    if (dl_out_mask_7) begin
      _T_5679 <= dl_out_data_7;
    end
    if (dl_out_mask_8) begin
      _T_5681 <= dl_out_data_8;
    end
    if (dl_out_mask_8) begin
      _T_5683 <= dl_out_data_8;
    end
    if (dl_out_mask_9) begin
      _T_5685 <= dl_out_data_9;
    end
    if (dl_out_mask_9) begin
      _T_5687 <= dl_out_data_9;
    end
    if (dl_out_mask_10) begin
      _T_5689 <= dl_out_data_10;
    end
    if (dl_out_mask_10) begin
      _T_5691 <= dl_out_data_10;
    end
    if (dl_out_mask_11) begin
      _T_5693 <= dl_out_data_11;
    end
    if (dl_out_mask_11) begin
      _T_5695 <= dl_out_data_11;
    end
    if (dl_out_mask_12) begin
      _T_5697 <= dl_out_data_12;
    end
    if (dl_out_mask_12) begin
      _T_5699 <= dl_out_data_12;
    end
    if (dl_out_mask_13) begin
      _T_5701 <= dl_out_data_13;
    end
    if (dl_out_mask_13) begin
      _T_5703 <= dl_out_data_13;
    end
    if (dl_out_mask_14) begin
      _T_5705 <= dl_out_data_14;
    end
    if (dl_out_mask_14) begin
      _T_5707 <= dl_out_data_14;
    end
    if (dl_out_mask_15) begin
      _T_5709 <= dl_out_data_15;
    end
    if (dl_out_mask_15) begin
      _T_5711 <= dl_out_data_15;
    end
    if (dl_out_mask_16) begin
      _T_5713 <= dl_out_data_16;
    end
    if (dl_out_mask_16) begin
      _T_5715 <= dl_out_data_16;
    end
    if (dl_out_mask_17) begin
      _T_5717 <= dl_out_data_17;
    end
    if (dl_out_mask_17) begin
      _T_5719 <= dl_out_data_17;
    end
    if (dl_out_mask_18) begin
      _T_5721 <= dl_out_data_18;
    end
    if (dl_out_mask_18) begin
      _T_5723 <= dl_out_data_18;
    end
    if (dl_out_mask_19) begin
      _T_5725 <= dl_out_data_19;
    end
    if (dl_out_mask_19) begin
      _T_5727 <= dl_out_data_19;
    end
    if (dl_out_mask_20) begin
      _T_5729 <= dl_out_data_20;
    end
    if (dl_out_mask_20) begin
      _T_5731 <= dl_out_data_20;
    end
    if (dl_out_mask_21) begin
      _T_5733 <= dl_out_data_21;
    end
    if (dl_out_mask_21) begin
      _T_5735 <= dl_out_data_21;
    end
    if (dl_out_mask_22) begin
      _T_5737 <= dl_out_data_22;
    end
    if (dl_out_mask_22) begin
      _T_5739 <= dl_out_data_22;
    end
    if (dl_out_mask_23) begin
      _T_5741 <= dl_out_data_23;
    end
    if (dl_out_mask_23) begin
      _T_5743 <= dl_out_data_23;
    end
    if (dl_out_mask_24) begin
      _T_5745 <= dl_out_data_24;
    end
    if (dl_out_mask_24) begin
      _T_5747 <= dl_out_data_24;
    end
    if (dl_out_mask_25) begin
      _T_5749 <= dl_out_data_25;
    end
    if (dl_out_mask_25) begin
      _T_5751 <= dl_out_data_25;
    end
    if (dl_out_mask_26) begin
      _T_5753 <= dl_out_data_26;
    end
    if (dl_out_mask_26) begin
      _T_5755 <= dl_out_data_26;
    end
    if (dl_out_mask_27) begin
      _T_5757 <= dl_out_data_27;
    end
    if (dl_out_mask_27) begin
      _T_5759 <= dl_out_data_27;
    end
    if (dl_out_mask_28) begin
      _T_5761 <= dl_out_data_28;
    end
    if (dl_out_mask_28) begin
      _T_5763 <= dl_out_data_28;
    end
    if (dl_out_mask_29) begin
      _T_5765 <= dl_out_data_29;
    end
    if (dl_out_mask_29) begin
      _T_5767 <= dl_out_data_29;
    end
    if (dl_out_mask_30) begin
      _T_5769 <= dl_out_data_30;
    end
    if (dl_out_mask_30) begin
      _T_5771 <= dl_out_data_30;
    end
    if (dl_out_mask_31) begin
      _T_5773 <= dl_out_data_31;
    end
    if (dl_out_mask_31) begin
      _T_5775 <= dl_out_data_31;
    end
    if (dl_out_mask_32) begin
      _T_5777 <= dl_out_data_32;
    end
    if (dl_out_mask_32) begin
      _T_5779 <= dl_out_data_32;
    end
    if (dl_out_mask_33) begin
      _T_5781 <= dl_out_data_33;
    end
    if (dl_out_mask_33) begin
      _T_5783 <= dl_out_data_33;
    end
    if (dl_out_mask_34) begin
      _T_5785 <= dl_out_data_34;
    end
    if (dl_out_mask_34) begin
      _T_5787 <= dl_out_data_34;
    end
    if (dl_out_mask_35) begin
      _T_5789 <= dl_out_data_35;
    end
    if (dl_out_mask_35) begin
      _T_5791 <= dl_out_data_35;
    end
    if (dl_out_mask_36) begin
      _T_5793 <= dl_out_data_36;
    end
    if (dl_out_mask_36) begin
      _T_5795 <= dl_out_data_36;
    end
    if (dl_out_mask_37) begin
      _T_5797 <= dl_out_data_37;
    end
    if (dl_out_mask_37) begin
      _T_5799 <= dl_out_data_37;
    end
    if (dl_out_mask_38) begin
      _T_5801 <= dl_out_data_38;
    end
    if (dl_out_mask_38) begin
      _T_5803 <= dl_out_data_38;
    end
    if (dl_out_mask_39) begin
      _T_5805 <= dl_out_data_39;
    end
    if (dl_out_mask_39) begin
      _T_5807 <= dl_out_data_39;
    end
    if (dl_out_mask_40) begin
      _T_5809 <= dl_out_data_40;
    end
    if (dl_out_mask_40) begin
      _T_5811 <= dl_out_data_40;
    end
    if (dl_out_mask_41) begin
      _T_5813 <= dl_out_data_41;
    end
    if (dl_out_mask_41) begin
      _T_5815 <= dl_out_data_41;
    end
    if (dl_out_mask_42) begin
      _T_5817 <= dl_out_data_42;
    end
    if (dl_out_mask_42) begin
      _T_5819 <= dl_out_data_42;
    end
    if (dl_out_mask_43) begin
      _T_5821 <= dl_out_data_43;
    end
    if (dl_out_mask_43) begin
      _T_5823 <= dl_out_data_43;
    end
    if (dl_out_mask_44) begin
      _T_5825 <= dl_out_data_44;
    end
    if (dl_out_mask_44) begin
      _T_5827 <= dl_out_data_44;
    end
    if (dl_out_mask_45) begin
      _T_5829 <= dl_out_data_45;
    end
    if (dl_out_mask_45) begin
      _T_5831 <= dl_out_data_45;
    end
    if (dl_out_mask_46) begin
      _T_5833 <= dl_out_data_46;
    end
    if (dl_out_mask_46) begin
      _T_5835 <= dl_out_data_46;
    end
    if (dl_out_mask_47) begin
      _T_5837 <= dl_out_data_47;
    end
    if (dl_out_mask_47) begin
      _T_5839 <= dl_out_data_47;
    end
    if (dl_out_mask_48) begin
      _T_5841 <= dl_out_data_48;
    end
    if (dl_out_mask_48) begin
      _T_5843 <= dl_out_data_48;
    end
    if (dl_out_mask_49) begin
      _T_5845 <= dl_out_data_49;
    end
    if (dl_out_mask_49) begin
      _T_5847 <= dl_out_data_49;
    end
    if (dl_out_mask_50) begin
      _T_5849 <= dl_out_data_50;
    end
    if (dl_out_mask_50) begin
      _T_5851 <= dl_out_data_50;
    end
    if (dl_out_mask_51) begin
      _T_5853 <= dl_out_data_51;
    end
    if (dl_out_mask_51) begin
      _T_5855 <= dl_out_data_51;
    end
    if (dl_out_mask_52) begin
      _T_5857 <= dl_out_data_52;
    end
    if (dl_out_mask_52) begin
      _T_5859 <= dl_out_data_52;
    end
    if (dl_out_mask_53) begin
      _T_5861 <= dl_out_data_53;
    end
    if (dl_out_mask_53) begin
      _T_5863 <= dl_out_data_53;
    end
    if (dl_out_mask_54) begin
      _T_5865 <= dl_out_data_54;
    end
    if (dl_out_mask_54) begin
      _T_5867 <= dl_out_data_54;
    end
    if (dl_out_mask_55) begin
      _T_5869 <= dl_out_data_55;
    end
    if (dl_out_mask_55) begin
      _T_5871 <= dl_out_data_55;
    end
    if (dl_out_mask_56) begin
      _T_5873 <= dl_out_data_56;
    end
    if (dl_out_mask_56) begin
      _T_5875 <= dl_out_data_56;
    end
    if (dl_out_mask_57) begin
      _T_5877 <= dl_out_data_57;
    end
    if (dl_out_mask_57) begin
      _T_5879 <= dl_out_data_57;
    end
    if (dl_out_mask_58) begin
      _T_5881 <= dl_out_data_58;
    end
    if (dl_out_mask_58) begin
      _T_5883 <= dl_out_data_58;
    end
    if (dl_out_mask_59) begin
      _T_5885 <= dl_out_data_59;
    end
    if (dl_out_mask_59) begin
      _T_5887 <= dl_out_data_59;
    end
    if (dl_out_mask_60) begin
      _T_5889 <= dl_out_data_60;
    end
    if (dl_out_mask_60) begin
      _T_5891 <= dl_out_data_60;
    end
    if (dl_out_mask_61) begin
      _T_5893 <= dl_out_data_61;
    end
    if (dl_out_mask_61) begin
      _T_5895 <= dl_out_data_61;
    end
    if (dl_out_mask_62) begin
      _T_5897 <= dl_out_data_62;
    end
    if (dl_out_mask_62) begin
      _T_5899 <= dl_out_data_62;
    end
    if (dl_out_mask_63) begin
      _T_5901 <= dl_out_data_63;
    end
    if (dl_out_mask_63) begin
      _T_5903 <= dl_out_data_63;
    end
  end
  always @(posedge io_nvdla_core_ng_clk) begin
    if (_T_207) begin
      dat_entry_st <= 15'h0;
    end else begin
      if (_T_638) begin
        if (io_sc2cdma_dat_pending_req) begin
          dat_entry_st <= 15'h0;
        end else begin
          if (is_dat_entry_st_wrap) begin
            dat_entry_st <= dat_entry_st_inc_wrap;
          end else begin
            dat_entry_st <= dat_entry_st_inc;
          end
        end
      end
    end
  end
endmodule
